
module my_DFF_1_0 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n3, n1, n2;

  DFFARX1 q_reg ( .D(n3), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n3) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_203 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X2 U2 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U3 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_202 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_201 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U2 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U3 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_200 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_199 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_198 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_197 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_nDFF_n8_0 ( clk, rst, e, d, q );
  input [7:0] d;
  output [7:0] q;
  input clk, rst, e;
  wire   n1;

  my_DFF_1_0 fx_0 ( .d(d[0]), .clk(clk), .rst(n1), .e(e), .q(q[0]) );
  my_DFF_1_203 fx_1 ( .d(d[1]), .clk(clk), .rst(n1), .e(e), .q(q[1]) );
  my_DFF_1_202 fx_2 ( .d(d[2]), .clk(clk), .rst(n1), .e(e), .q(q[2]) );
  my_DFF_1_201 fx_3 ( .d(d[3]), .clk(clk), .rst(n1), .e(e), .q(q[3]) );
  my_DFF_1_200 fx_4 ( .d(d[4]), .clk(clk), .rst(n1), .e(e), .q(q[4]) );
  my_DFF_1_199 fx_5 ( .d(d[5]), .clk(clk), .rst(n1), .e(e), .q(q[5]) );
  my_DFF_1_198 fx_6 ( .d(d[6]), .clk(clk), .rst(n1), .e(e), .q(q[6]) );
  my_DFF_1_197 fx_7 ( .d(d[7]), .clk(clk), .rst(n1), .e(e), .q(q[7]) );
  NBUFFX2 U1 ( .IN(rst), .Q(n1) );
endmodule


module inst_ram_1 ( clk, R, address, dataout, MFC );
  input [7:0] address;
  output [7:0] dataout;
  input clk, R;
  output MFC;

  assign dataout[7] = 1'b0;
  assign dataout[6] = 1'b0;
  assign dataout[5] = 1'b0;
  assign dataout[4] = 1'b0;
  assign dataout[3] = 1'b0;
  assign dataout[2] = 1'b0;
  assign dataout[1] = 1'b0;
  assign dataout[0] = 1'b0;

  DFFNX1 MFC_reg ( .D(R), .CLK(clk), .Q(MFC) );
endmodule


module my_DFF_1_196 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_195 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_194 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_193 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_192 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_191 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_190 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_189 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_188 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_187 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_186 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_185 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_184 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_183 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_182 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_181 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_180 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_179 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_178 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_177 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_176 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_175 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_174 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_173 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_172 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_171 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_170 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_169 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_168 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_167 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_166 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_165 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_nDFF_n32_0 ( clk, rst, e, d, q );
  input [31:0] d;
  output [31:0] q;
  input clk, rst, e;
  wire   n1, n2, n3;

  my_DFF_1_196 fx_0 ( .d(d[0]), .clk(clk), .rst(rst), .e(n3), .q(q[0]) );
  my_DFF_1_195 fx_1 ( .d(d[1]), .clk(clk), .rst(rst), .e(n3), .q(q[1]) );
  my_DFF_1_194 fx_2 ( .d(d[2]), .clk(clk), .rst(rst), .e(n3), .q(q[2]) );
  my_DFF_1_193 fx_3 ( .d(d[3]), .clk(clk), .rst(rst), .e(n3), .q(q[3]) );
  my_DFF_1_192 fx_4 ( .d(d[4]), .clk(clk), .rst(rst), .e(n3), .q(q[4]) );
  my_DFF_1_191 fx_5 ( .d(d[5]), .clk(clk), .rst(rst), .e(n3), .q(q[5]) );
  my_DFF_1_190 fx_6 ( .d(d[6]), .clk(clk), .rst(rst), .e(n3), .q(q[6]) );
  my_DFF_1_189 fx_7 ( .d(d[7]), .clk(clk), .rst(rst), .e(n3), .q(q[7]) );
  my_DFF_1_188 fx_8 ( .d(d[8]), .clk(clk), .rst(rst), .e(n2), .q(q[8]) );
  my_DFF_1_187 fx_9 ( .d(d[9]), .clk(clk), .rst(rst), .e(n2), .q(q[9]) );
  my_DFF_1_186 fx_10 ( .d(d[10]), .clk(clk), .rst(rst), .e(n2), .q(q[10]) );
  my_DFF_1_185 fx_11 ( .d(d[11]), .clk(clk), .rst(rst), .e(n2), .q(q[11]) );
  my_DFF_1_184 fx_12 ( .d(d[12]), .clk(clk), .rst(rst), .e(n2), .q(q[12]) );
  my_DFF_1_183 fx_13 ( .d(d[13]), .clk(clk), .rst(rst), .e(n2), .q(q[13]) );
  my_DFF_1_182 fx_14 ( .d(d[14]), .clk(clk), .rst(rst), .e(n2), .q(q[14]) );
  my_DFF_1_181 fx_15 ( .d(d[15]), .clk(clk), .rst(rst), .e(n2), .q(q[15]) );
  my_DFF_1_180 fx_16 ( .d(d[16]), .clk(clk), .rst(rst), .e(n2), .q(q[16]) );
  my_DFF_1_179 fx_17 ( .d(d[17]), .clk(clk), .rst(rst), .e(n2), .q(q[17]) );
  my_DFF_1_178 fx_18 ( .d(d[18]), .clk(clk), .rst(rst), .e(n2), .q(q[18]) );
  my_DFF_1_177 fx_19 ( .d(d[19]), .clk(clk), .rst(rst), .e(n2), .q(q[19]) );
  my_DFF_1_176 fx_20 ( .d(d[20]), .clk(clk), .rst(rst), .e(n1), .q(q[20]) );
  my_DFF_1_175 fx_21 ( .d(d[21]), .clk(clk), .rst(rst), .e(n1), .q(q[21]) );
  my_DFF_1_174 fx_22 ( .d(d[22]), .clk(clk), .rst(rst), .e(n1), .q(q[22]) );
  my_DFF_1_173 fx_23 ( .d(d[23]), .clk(clk), .rst(rst), .e(n1), .q(q[23]) );
  my_DFF_1_172 fx_24 ( .d(d[24]), .clk(clk), .rst(rst), .e(n1), .q(q[24]) );
  my_DFF_1_171 fx_25 ( .d(d[25]), .clk(clk), .rst(rst), .e(n1), .q(q[25]) );
  my_DFF_1_170 fx_26 ( .d(d[26]), .clk(clk), .rst(rst), .e(n1), .q(q[26]) );
  my_DFF_1_169 fx_27 ( .d(d[27]), .clk(clk), .rst(rst), .e(n1), .q(q[27]) );
  my_DFF_1_168 fx_28 ( .d(d[28]), .clk(clk), .rst(rst), .e(n1), .q(q[28]) );
  my_DFF_1_167 fx_29 ( .d(d[29]), .clk(clk), .rst(rst), .e(n1), .q(q[29]) );
  my_DFF_1_166 fx_30 ( .d(d[30]), .clk(clk), .rst(rst), .e(n1), .q(q[30]) );
  my_DFF_1_165 fx_31 ( .d(d[31]), .clk(clk), .rst(rst), .e(n1), .q(q[31]) );
  NBUFFX2 U1 ( .IN(e), .Q(n2) );
  NBUFFX2 U2 ( .IN(e), .Q(n1) );
  NBUFFX2 U3 ( .IN(e), .Q(n3) );
endmodule


module CU_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[7]), .IN2(A[7]), .Q(SUM[7]) );
endmodule


module CU ( clk, rst, INT_IN, stall, ret_Ex, ret_Mem, ret_WB, branch, EX_RTI, 
        ret_PC, target_address, IF_ID, reg_R, inst_R, stall_en, IR_rst, f1_en, 
        f2_en, imm_en, Rs1, Rs2, Rd, acc_mode, NOP, offset_en, offset, alu_op, 
        change_flags, branch_mode, ret, PC_src, push_PC, push_flags, 
        return_address, return_address_src, flags_src, pre_RTI, pre_pop_flags, 
        PCin );
  input [7:0] ret_PC;
  input [7:0] target_address;
  input [31:0] IF_ID;
  output [1:0] Rs1;
  output [1:0] Rs2;
  output [1:0] Rd;
  output [2:0] acc_mode;
  output [7:0] offset;
  output [3:0] alu_op;
  output [2:0] branch_mode;
  output [7:0] return_address;
  output [7:0] PCin;
  input clk, rst, INT_IN, stall, ret_Ex, ret_Mem, ret_WB, branch, EX_RTI;
  output reg_R, inst_R, stall_en, IR_rst, f1_en, f2_en, imm_en, NOP, offset_en,
         change_flags, ret, PC_src, push_PC, push_flags, return_address_src,
         flags_src, pre_RTI, pre_pop_flags;
  wire   EX_RTI, \IF_ID[1] , \IF_ID[0] , INT, N37, used_INT, N57, N59, N60,
         N61, N62, N63, N64, N65, N66, N92, N93, N94, N95, N96, N97, N98, N99,
         N122, N135, N144, N476, N493, N690, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n30, n31, n32, n33, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, inst_R, n156, n157, n158;
  assign reg_R = 1'b1;
  assign offset[1] = 1'b0;
  assign offset[2] = 1'b0;
  assign offset[3] = 1'b0;
  assign offset[4] = 1'b0;
  assign offset[5] = 1'b0;
  assign offset[6] = 1'b0;
  assign offset[7] = 1'b0;
  assign pre_pop_flags = EX_RTI;
  assign return_address_src = IF_ID[17];
  assign flags_src = IF_ID[16];
  assign push_PC = IF_ID[16];
  assign Rs2[1] = \IF_ID[1] ;
  assign \IF_ID[1]  = IF_ID[1];
  assign Rs2[0] = \IF_ID[0] ;
  assign \IF_ID[0]  = IF_ID[0];
  assign push_flags = INT;
  assign pre_RTI = N122;
  assign IR_rst = N135;
  assign ret = N144;
  assign offset_en = N476;
  assign offset[0] = N493;
  assign change_flags = N690;
  assign stall_en = inst_R;

  DFFARX1 INT_reg ( .D(1'b1), .CLK(used_INT), .RSTB(n158), .Q(INT) );
  OR2X1 U97 ( .IN1(n34), .IN2(INT_IN), .Q(used_INT) );
  AO22X1 U98 ( .IN1(N99), .IN2(INT), .IN3(IF_ID[25]), .IN4(n38), .Q(
        return_address[7]) );
  AO22X1 U99 ( .IN1(N98), .IN2(INT), .IN3(IF_ID[24]), .IN4(n38), .Q(
        return_address[6]) );
  AO22X1 U100 ( .IN1(N97), .IN2(INT), .IN3(IF_ID[23]), .IN4(n38), .Q(
        return_address[5]) );
  AO22X1 U101 ( .IN1(N96), .IN2(INT), .IN3(IF_ID[22]), .IN4(n38), .Q(
        return_address[4]) );
  AO22X1 U102 ( .IN1(N95), .IN2(INT), .IN3(IF_ID[21]), .IN4(n38), .Q(
        return_address[3]) );
  AO22X1 U103 ( .IN1(N94), .IN2(INT), .IN3(IF_ID[20]), .IN4(n38), .Q(
        return_address[2]) );
  AO22X1 U104 ( .IN1(N93), .IN2(INT), .IN3(IF_ID[19]), .IN4(n38), .Q(
        return_address[1]) );
  AO22X1 U105 ( .IN1(N92), .IN2(INT), .IN3(IF_ID[18]), .IN4(n38), .Q(
        return_address[0]) );
  AND3X1 U106 ( .IN1(n40), .IN2(n156), .IN3(n39), .Q(f2_en) );
  NAND4X0 U107 ( .IN1(n41), .IN2(n42), .IN3(n43), .IN4(n44), .QN(n40) );
  OA21X1 U108 ( .IN1(n19), .IN2(n45), .IN3(n46), .Q(n44) );
  XNOR2X1 U109 ( .IN1(n37), .IN2(n151), .Q(n46) );
  NAND3X0 U110 ( .IN1(n153), .IN2(n49), .IN3(n18), .QN(n47) );
  NAND3X0 U111 ( .IN1(n50), .IN2(n51), .IN3(n52), .QN(n49) );
  NAND4X0 U112 ( .IN1(n18), .IN2(n50), .IN3(n51), .IN4(n53), .QN(n42) );
  NAND3X0 U113 ( .IN1(n153), .IN2(n54), .IN3(n55), .QN(n41) );
  AO221X1 U114 ( .IN1(n19), .IN2(n56), .IN3(n57), .IN4(n53), .IN5(n58), .Q(
        f1_en) );
  NAND3X0 U115 ( .IN1(n153), .IN2(n54), .IN3(n149), .QN(n59) );
  NAND3X0 U116 ( .IN1(n51), .IN2(n53), .IN3(n52), .QN(n45) );
  NAND3X0 U117 ( .IN1(n61), .IN2(n62), .IN3(n63), .QN(branch_mode[2]) );
  NAND3X0 U118 ( .IN1(n65), .IN2(n66), .IN3(n63), .QN(branch_mode[1]) );
  NAND4X0 U119 ( .IN1(n67), .IN2(n66), .IN3(n62), .IN4(n68), .QN(
        branch_mode[0]) );
  AND2X1 U120 ( .IN1(n69), .IN2(n19), .Q(n64) );
  OA21X1 U121 ( .IN1(n147), .IN2(n27), .IN3(n24), .Q(alu_op[3]) );
  AND4X1 U122 ( .IN1(n73), .IN2(n74), .IN3(n75), .IN4(n76), .Q(n71) );
  NAND3X0 U123 ( .IN1(n82), .IN2(n83), .IN3(n73), .QN(n79) );
  AO21X1 U124 ( .IN1(n24), .IN2(n84), .IN3(n78), .Q(alu_op[0]) );
  NAND3X0 U125 ( .IN1(n19), .IN2(n48), .IN3(n150), .QN(n86) );
  NAND4X0 U126 ( .IN1(n87), .IN2(n83), .IN3(n73), .IN4(n88), .QN(n84) );
  OA221X1 U127 ( .IN1(n51), .IN2(n143), .IN3(n36), .IN4(n75), .IN5(n146), .Q(
        n88) );
  NAND3X0 U128 ( .IN1(n91), .IN2(n92), .IN3(n93), .QN(n72) );
  AO21X1 U129 ( .IN1(n35), .IN2(n89), .IN3(n18), .Q(n91) );
  NAND4X0 U130 ( .IN1(n25), .IN2(n76), .IN3(n94), .IN4(n85), .QN(acc_mode[2])
         );
  NAND3X0 U131 ( .IN1(n76), .IN2(n94), .IN3(n95), .QN(acc_mode[1]) );
  NAND3X0 U132 ( .IN1(n96), .IN2(n85), .IN3(n25), .QN(n95) );
  NAND3X0 U133 ( .IN1(n99), .IN2(n36), .IN3(n151), .QN(n98) );
  AO21X1 U134 ( .IN1(n94), .IN2(n100), .IN3(n27), .Q(acc_mode[0]) );
  OA22X1 U135 ( .IN1(n143), .IN2(n52), .IN3(n143), .IN4(n51), .Q(n76) );
  OAI21X1 U136 ( .IN1(n102), .IN2(n103), .IN3(n85), .QN(n100) );
  OA21X1 U137 ( .IN1(n55), .IN2(n92), .IN3(n97), .Q(n102) );
  AND2X1 U138 ( .IN1(n25), .IN2(n97), .Q(n93) );
  AND2X1 U139 ( .IN1(n105), .IN2(n106), .Q(n97) );
  AO22X1 U140 ( .IN1(IF_ID[3]), .IN2(n108), .IN3(\IF_ID[1] ), .IN4(n109), .Q(
        Rd[1]) );
  AO22X1 U141 ( .IN1(IF_ID[2]), .IN2(n108), .IN3(\IF_ID[0] ), .IN4(n109), .Q(
        Rd[0]) );
  NAND3X0 U142 ( .IN1(n92), .IN2(n101), .IN3(n110), .QN(n109) );
  AO21X1 U143 ( .IN1(n153), .IN2(n37), .IN3(n148), .Q(n111) );
  AO22X1 U144 ( .IN1(n57), .IN2(n53), .IN3(n112), .IN4(n36), .Q(n108) );
  AO221X1 U145 ( .IN1(N66), .IN2(n113), .IN3(ret_PC[7]), .IN4(n114), .IN5(n115), .Q(PCin[7]) );
  AO221X1 U147 ( .IN1(N65), .IN2(n113), .IN3(ret_PC[6]), .IN4(n114), .IN5(n117), .Q(PCin[6]) );
  AO22X1 U148 ( .IN1(n154), .IN2(IF_ID[6]), .IN3(target_address[6]), .IN4(n5), 
        .Q(n117) );
  AO221X1 U149 ( .IN1(N64), .IN2(n113), .IN3(ret_PC[5]), .IN4(n114), .IN5(n118), .Q(PCin[5]) );
  AO221X1 U151 ( .IN1(N63), .IN2(n113), .IN3(ret_PC[4]), .IN4(n114), .IN5(n119), .Q(PCin[4]) );
  AO22X1 U152 ( .IN1(n154), .IN2(IF_ID[4]), .IN3(target_address[4]), .IN4(n5), 
        .Q(n119) );
  AO221X1 U153 ( .IN1(N62), .IN2(n113), .IN3(ret_PC[3]), .IN4(n114), .IN5(n120), .Q(PCin[3]) );
  AO22X1 U154 ( .IN1(n154), .IN2(IF_ID[3]), .IN3(target_address[3]), .IN4(n116), .Q(n120) );
  AO221X1 U155 ( .IN1(N61), .IN2(n113), .IN3(ret_PC[2]), .IN4(n114), .IN5(n121), .Q(PCin[2]) );
  AO22X1 U156 ( .IN1(n154), .IN2(IF_ID[2]), .IN3(target_address[2]), .IN4(n116), .Q(n121) );
  AO221X1 U157 ( .IN1(N60), .IN2(n113), .IN3(ret_PC[1]), .IN4(n114), .IN5(n122), .Q(PCin[1]) );
  AO22X1 U163 ( .IN1(n154), .IN2(\IF_ID[0] ), .IN3(n127), .IN4(n128), .Q(
        PCin[0]) );
  AO221X1 U164 ( .IN1(n129), .IN2(n124), .IN3(target_address[0]), .IN4(n6), 
        .IN5(n123), .Q(n127) );
  AO22X1 U166 ( .IN1(ret_PC[0]), .IN2(n157), .IN3(N59), .IN4(n126), .Q(n129)
         );
  NAND3X0 U167 ( .IN1(n130), .IN2(n156), .IN3(n39), .QN(NOP) );
  NAND3X0 U168 ( .IN1(n21), .IN2(n20), .IN3(n131), .QN(n130) );
  AO221X1 U169 ( .IN1(n112), .IN2(n54), .IN3(n132), .IN4(n36), .IN5(n133), .Q(
        n131) );
  AO22X1 U170 ( .IN1(n152), .IN2(n37), .IN3(n18), .IN4(n53), .Q(n133) );
  NAND4X0 U171 ( .IN1(n134), .IN2(n135), .IN3(n90), .IN4(n89), .QN(N690) );
  AND3X1 U172 ( .IN1(n37), .IN2(n48), .IN3(n153), .Q(n69) );
  NAND3X0 U173 ( .IN1(n36), .IN2(n53), .IN3(n152), .QN(n135) );
  OAI21X1 U174 ( .IN1(IF_ID[17]), .IN2(stall), .IN3(n20), .QN(N57) );
  NAND4X0 U175 ( .IN1(n136), .IN2(n107), .IN3(n138), .IN4(n139), .QN(N476) );
  AND2X1 U176 ( .IN1(n60), .IN2(n92), .Q(n138) );
  NAND3X0 U177 ( .IN1(n153), .IN2(n36), .IN3(n149), .QN(n60) );
  OA21X1 U178 ( .IN1(n145), .IN2(n54), .IN3(n39), .Q(n107) );
  AOI21X1 U179 ( .IN1(n137), .IN2(n140), .IN3(n31), .QN(n136) );
  OA21X1 U180 ( .IN1(n145), .IN2(n50), .IN3(n156), .Q(n106) );
  AO21X1 U181 ( .IN1(clk), .IN2(INT), .IN3(rst), .Q(N37) );
  OAI21X1 U182 ( .IN1(rst), .IN2(n142), .IN3(n128), .QN(N135) );
  AND2X1 U183 ( .IN1(n70), .IN2(n26), .Q(n141) );
  AND2X1 U184 ( .IN1(n70), .IN2(n32), .Q(N122) );
  AND2X1 U185 ( .IN1(n137), .IN2(n18), .Q(n70) );
  AND2X1 U186 ( .IN1(n112), .IN2(n153), .Q(n137) );
  CU_DW01_inc_0 add_85 ( .A(IF_ID[15:8]), .SUM({N99, N98, N97, N96, N95, N94, 
        N93, N92}) );
  DELLN1X2 U3 ( .IN(branch), .Q(n2) );
  AND2X1 U4 ( .IN1(branch), .IN2(n20), .Q(n6) );
  AO22X1 U5 ( .IN1(n154), .IN2(IF_ID[5]), .IN3(target_address[5]), .IN4(n116), 
        .Q(n118) );
  INVX0 U6 ( .IN(n2), .QN(n21) );
  NOR2X0 U7 ( .IN1(n6), .IN2(n9), .QN(n1) );
  NAND2X0 U8 ( .IN1(n154), .IN2(\IF_ID[1] ), .QN(n3) );
  NAND2X0 U9 ( .IN1(target_address[1]), .IN2(n5), .QN(n4) );
  NAND2X0 U10 ( .IN1(n3), .IN2(n4), .QN(n122) );
  NAND2X0 U11 ( .IN1(branch), .IN2(n20), .QN(n124) );
  NOR2X0 U12 ( .IN1(n124), .IN2(n8), .QN(n5) );
  NOR2X0 U13 ( .IN1(n124), .IN2(n8), .QN(n116) );
  INVX0 U14 ( .IN(n7), .QN(n8) );
  AND2X1 U15 ( .IN1(INT), .IN2(n20), .Q(n123) );
  NOR2X0 U16 ( .IN1(n154), .IN2(n123), .QN(n7) );
  AO22X1 U17 ( .IN1(n154), .IN2(IF_ID[7]), .IN3(target_address[7]), .IN4(n5), 
        .Q(n115) );
  OR2X1 U18 ( .IN1(n154), .IN2(n123), .Q(n9) );
  NOR2X0 U19 ( .IN1(n6), .IN2(n9), .QN(n125) );
  INVX0 U20 ( .IN(n74), .QN(n22) );
  NOR2X0 U21 ( .IN1(N122), .IN2(n141), .QN(n105) );
  INVX0 U22 ( .IN(n72), .QN(n24) );
  INVX0 U23 ( .IN(n57), .QN(n148) );
  INVX0 U24 ( .IN(n103), .QN(n25) );
  INVX0 U25 ( .IN(n35), .QN(n151) );
  INVX0 U26 ( .IN(n68), .QN(PC_src) );
  INVX0 U27 ( .IN(n81), .QN(n143) );
  NAND2X0 U28 ( .IN1(n81), .IN2(n23), .QN(n74) );
  NAND2X0 U29 ( .IN1(n150), .IN2(n17), .QN(n134) );
  AND2X1 U30 ( .IN1(n157), .IN2(n1), .Q(n114) );
  NAND2X0 U31 ( .IN1(n70), .IN2(n30), .QN(n68) );
  NAND2X0 U32 ( .IN1(n149), .IN2(n152), .QN(n57) );
  NAND2X0 U33 ( .IN1(n107), .IN2(n68), .QN(n103) );
  INVX0 U34 ( .IN(n104), .QN(n145) );
  NBUFFX2 U35 ( .IN(n144), .Q(n18) );
  NOR2X0 U36 ( .IN1(n101), .IN2(n17), .QN(n81) );
  INVX0 U37 ( .IN(n90), .QN(n147) );
  NAND2X0 U38 ( .IN1(n147), .IN2(n26), .QN(n82) );
  NAND2X0 U39 ( .IN1(n153), .IN2(n152), .QN(n35) );
  INVX0 U40 ( .IN(n132), .QN(n150) );
  NOR2X0 U41 ( .IN1(n19), .IN2(n30), .QN(n55) );
  NOR2X0 U42 ( .IN1(n92), .IN2(n17), .QN(imm_en) );
  NAND2X0 U43 ( .IN1(n104), .IN2(n26), .QN(n85) );
  NAND2X0 U44 ( .IN1(n81), .IN2(n30), .QN(n73) );
  NAND2X0 U45 ( .IN1(n32), .IN2(n64), .QN(n62) );
  NAND2X0 U46 ( .IN1(n30), .IN2(n64), .QN(n66) );
  NAND2X0 U47 ( .IN1(n104), .IN2(n32), .QN(n94) );
  NAND2X0 U48 ( .IN1(n147), .IN2(n32), .QN(n83) );
  NAND2X0 U49 ( .IN1(n150), .IN2(n152), .QN(n75) );
  NAND2X0 U50 ( .IN1(n63), .IN2(n89), .QN(n80) );
  NAND2X0 U51 ( .IN1(n147), .IN2(n30), .QN(n87) );
  NAND2X0 U52 ( .IN1(n35), .IN2(n45), .QN(n56) );
  INVX0 U53 ( .IN(n76), .QN(n27) );
  NBUFFX2 U54 ( .IN(n144), .Q(n17) );
  NBUFFX2 U55 ( .IN(n144), .Q(n19) );
  INVX0 U56 ( .IN(n54), .QN(n23) );
  INVX0 U57 ( .IN(rst), .QN(n20) );
  INVX0 U58 ( .IN(stall), .QN(inst_R) );
  INVX0 U59 ( .IN(n48), .QN(n152) );
  INVX0 U60 ( .IN(n53), .QN(n153) );
  NOR2X0 U61 ( .IN1(n101), .IN2(n36), .QN(n104) );
  INVX0 U62 ( .IN(n52), .QN(n26) );
  NOR2X0 U63 ( .IN1(n37), .IN2(n152), .QN(n112) );
  NAND2X0 U64 ( .IN1(n148), .IN2(n53), .QN(n101) );
  INVX0 U65 ( .IN(n37), .QN(n149) );
  NAND2X0 U66 ( .IN1(n93), .IN2(n28), .QN(Rs1[0]) );
  NAND2X0 U67 ( .IN1(n93), .IN2(n33), .QN(Rs1[1]) );
  INVX0 U68 ( .IN(n36), .QN(n144) );
  INVX0 U69 ( .IN(n50), .QN(n30) );
  NAND2X0 U70 ( .IN1(n47), .IN2(n48), .QN(n43) );
  INVX0 U71 ( .IN(n128), .QN(n154) );
  NAND2X0 U72 ( .IN1(n111), .IN2(n36), .QN(n110) );
  INVX0 U73 ( .IN(n51), .QN(n32) );
  NAND2X0 U74 ( .IN1(n137), .IN2(n36), .QN(n63) );
  INVX0 U75 ( .IN(n80), .QN(n146) );
  NAND2X0 U76 ( .IN1(n151), .IN2(n37), .QN(n92) );
  NAND2X0 U77 ( .IN1(n112), .IN2(n53), .QN(n89) );
  NAND2X0 U78 ( .IN1(n33), .IN2(n28), .QN(n54) );
  NAND2X0 U79 ( .IN1(n69), .IN2(n36), .QN(n90) );
  NAND2X0 U80 ( .IN1(n51), .IN2(n52), .QN(n140) );
  INVX0 U81 ( .IN(n106), .QN(n31) );
  NAND2X0 U82 ( .IN1(n53), .IN2(n37), .QN(n132) );
  NAND2X0 U83 ( .IN1(n85), .IN2(n86), .QN(n78) );
  NAND2X0 U84 ( .IN1(n97), .IN2(n98), .QN(n96) );
  NAND2X0 U85 ( .IN1(n37), .IN2(n52), .QN(n99) );
  INVX0 U86 ( .IN(n126), .QN(n157) );
  XNOR2X1 U87 ( .IN1(n16), .IN2(IF_ID[15]), .Q(N66) );
  AND2X1 U88 ( .IN1(N57), .IN2(IF_ID[8]), .Q(n10) );
  AND2X1 U89 ( .IN1(n10), .IN2(IF_ID[9]), .Q(n11) );
  AND2X1 U90 ( .IN1(n11), .IN2(IF_ID[10]), .Q(n12) );
  AND2X1 U91 ( .IN1(n12), .IN2(IF_ID[11]), .Q(n13) );
  AND2X1 U92 ( .IN1(n13), .IN2(IF_ID[12]), .Q(n14) );
  AND2X1 U93 ( .IN1(n14), .IN2(IF_ID[13]), .Q(n15) );
  NAND2X0 U94 ( .IN1(n15), .IN2(IF_ID[14]), .QN(n16) );
  NOR2X0 U95 ( .IN1(IF_ID[17]), .IN2(IF_ID[16]), .QN(n39) );
  NAND2X0 U96 ( .IN1(IF_ID[4]), .IN2(n39), .QN(n36) );
  NAND2X0 U146 ( .IN1(IF_ID[5]), .IN2(n39), .QN(n37) );
  NAND2X0 U150 ( .IN1(IF_ID[7]), .IN2(n39), .QN(n53) );
  NAND2X0 U158 ( .IN1(IF_ID[3]), .IN2(n28), .QN(n52) );
  INVX0 U159 ( .IN(IF_ID[2]), .QN(n28) );
  NAND2X0 U160 ( .IN1(IF_ID[6]), .IN2(n39), .QN(n48) );
  NOR2X0 U161 ( .IN1(n71), .IN2(n72), .QN(alu_op[2]) );
  NOR2X0 U162 ( .IN1(n77), .IN2(n78), .QN(alu_op[1]) );
  NOR4X0 U165 ( .IN1(n79), .IN2(n80), .IN3(n22), .IN4(n72), .QN(n77) );
  NAND2X0 U187 ( .IN1(IF_ID[3]), .IN2(IF_ID[2]), .QN(n51) );
  INVX0 U188 ( .IN(IF_ID[3]), .QN(n33) );
  NAND2X0 U189 ( .IN1(IF_ID[2]), .IN2(n33), .QN(n50) );
  NOR2X0 U190 ( .IN1(rst), .IN2(n105), .QN(N144) );
  NAND2X0 U191 ( .IN1(n136), .IN2(n63), .QN(N493) );
  NAND2X0 U192 ( .IN1(n23), .IN2(n64), .QN(n65) );
  NAND2X0 U193 ( .IN1(n26), .IN2(n64), .QN(n61) );
  NAND2X0 U194 ( .IN1(n30), .IN2(n137), .QN(n139) );
  NAND2X0 U195 ( .IN1(n59), .IN2(n60), .QN(n58) );
  NAND2X0 U196 ( .IN1(n70), .IN2(n23), .QN(n67) );
  NAND2X0 U197 ( .IN1(ret_WB), .IN2(n20), .QN(n126) );
  NAND2X0 U198 ( .IN1(IF_ID[16]), .IN2(n20), .QN(n128) );
  INVX0 U199 ( .IN(EX_RTI), .QN(n156) );
  NOR2X0 U200 ( .IN1(n39), .IN2(INT), .QN(n38) );
  INVX0 U201 ( .IN(N37), .QN(n158) );
  NOR4X0 U202 ( .IN1(ret_Mem), .IN2(ret_Ex), .IN3(imm_en), .IN4(n141), .QN(
        n142) );
  NOR4X0 U203 ( .IN1(rst), .IN2(n35), .IN3(n36), .IN4(n37), .QN(n34) );
  XOR2X1 U204 ( .IN1(N57), .IN2(IF_ID[8]), .Q(N59) );
  XOR2X1 U205 ( .IN1(n10), .IN2(IF_ID[9]), .Q(N60) );
  XOR2X1 U206 ( .IN1(n11), .IN2(IF_ID[10]), .Q(N61) );
  XOR2X1 U207 ( .IN1(n12), .IN2(IF_ID[11]), .Q(N62) );
  XOR2X1 U208 ( .IN1(n13), .IN2(IF_ID[12]), .Q(N63) );
  XOR2X1 U209 ( .IN1(n14), .IN2(IF_ID[13]), .Q(N64) );
  XOR2X1 U210 ( .IN1(n15), .IN2(IF_ID[14]), .Q(N65) );
  AND2X2 U211 ( .IN1(n125), .IN2(n126), .Q(n113) );
endmodule


module my_DFF_1_32 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_31 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_30 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_29 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_28 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_27 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_26 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_25 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_nDFF_n8_4 ( clk, rst, e, d, q );
  input [7:0] d;
  output [7:0] q;
  input clk, rst, e;
  wire   n1;

  my_DFF_1_32 fx_0 ( .d(d[0]), .clk(clk), .rst(n1), .e(e), .q(q[0]) );
  my_DFF_1_31 fx_1 ( .d(d[1]), .clk(clk), .rst(n1), .e(e), .q(q[1]) );
  my_DFF_1_30 fx_2 ( .d(d[2]), .clk(clk), .rst(n1), .e(e), .q(q[2]) );
  my_DFF_1_29 fx_3 ( .d(d[3]), .clk(clk), .rst(n1), .e(e), .q(q[3]) );
  my_DFF_1_28 fx_4 ( .d(d[4]), .clk(clk), .rst(n1), .e(e), .q(q[4]) );
  my_DFF_1_27 fx_5 ( .d(d[5]), .clk(clk), .rst(n1), .e(e), .q(q[5]) );
  my_DFF_1_26 fx_6 ( .d(d[6]), .clk(clk), .rst(n1), .e(e), .q(q[6]) );
  my_DFF_1_25 fx_7 ( .d(d[7]), .clk(clk), .rst(n1), .e(e), .q(q[7]) );
  NBUFFX2 U1 ( .IN(rst), .Q(n1) );
endmodule


module my_DFF_1_24 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_23 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_22 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_21 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_20 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_19 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_18 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_17 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_nDFF_n8_3 ( clk, rst, e, d, q );
  input [7:0] d;
  output [7:0] q;
  input clk, rst, e;
  wire   n1;

  my_DFF_1_24 fx_0 ( .d(d[0]), .clk(clk), .rst(n1), .e(e), .q(q[0]) );
  my_DFF_1_23 fx_1 ( .d(d[1]), .clk(clk), .rst(n1), .e(e), .q(q[1]) );
  my_DFF_1_22 fx_2 ( .d(d[2]), .clk(clk), .rst(n1), .e(e), .q(q[2]) );
  my_DFF_1_21 fx_3 ( .d(d[3]), .clk(clk), .rst(n1), .e(e), .q(q[3]) );
  my_DFF_1_20 fx_4 ( .d(d[4]), .clk(clk), .rst(n1), .e(e), .q(q[4]) );
  my_DFF_1_19 fx_5 ( .d(d[5]), .clk(clk), .rst(n1), .e(e), .q(q[5]) );
  my_DFF_1_18 fx_6 ( .d(d[6]), .clk(clk), .rst(n1), .e(e), .q(q[6]) );
  my_DFF_1_17 fx_7 ( .d(d[7]), .clk(clk), .rst(n1), .e(e), .q(q[7]) );
  NBUFFX2 U1 ( .IN(rst), .Q(n1) );
endmodule


module my_DFF_1_16 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_15 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_14 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_13 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_12 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_11 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_10 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_9 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_nDFF_n8_2 ( clk, rst, e, d, q );
  input [7:0] d;
  output [7:0] q;
  input clk, rst, e;
  wire   n1;

  my_DFF_1_16 fx_0 ( .d(d[0]), .clk(clk), .rst(n1), .e(e), .q(q[0]) );
  my_DFF_1_15 fx_1 ( .d(d[1]), .clk(clk), .rst(n1), .e(e), .q(q[1]) );
  my_DFF_1_14 fx_2 ( .d(d[2]), .clk(clk), .rst(n1), .e(e), .q(q[2]) );
  my_DFF_1_13 fx_3 ( .d(d[3]), .clk(clk), .rst(n1), .e(e), .q(q[3]) );
  my_DFF_1_12 fx_4 ( .d(d[4]), .clk(clk), .rst(n1), .e(e), .q(q[4]) );
  my_DFF_1_11 fx_5 ( .d(d[5]), .clk(clk), .rst(n1), .e(e), .q(q[5]) );
  my_DFF_1_10 fx_6 ( .d(d[6]), .clk(clk), .rst(n1), .e(e), .q(q[6]) );
  my_DFF_1_9 fx_7 ( .d(d[7]), .clk(clk), .rst(n1), .e(e), .q(q[7]) );
  NBUFFX2 U1 ( .IN(rst), .Q(n1) );
endmodule


module my_DFF_1_8 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_7 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_6 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_5 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_4 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_3 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_2 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_DFF_1_1 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(e), .QN(n1) );
  INVX0 U4 ( .IN(rst), .QN(n2) );
endmodule


module my_nDFF_n8_1 ( clk, rst, e, d, q );
  input [7:0] d;
  output [7:0] q;
  input clk, rst, e;


  my_DFF_1_8 fx_0 ( .d(d[0]), .clk(clk), .rst(rst), .e(e), .q(q[0]) );
  my_DFF_1_7 fx_1 ( .d(d[1]), .clk(clk), .rst(rst), .e(e), .q(q[1]) );
  my_DFF_1_6 fx_2 ( .d(d[2]), .clk(clk), .rst(rst), .e(e), .q(q[2]) );
  my_DFF_1_5 fx_3 ( .d(d[3]), .clk(clk), .rst(rst), .e(e), .q(q[3]) );
  my_DFF_1_4 fx_4 ( .d(d[4]), .clk(clk), .rst(rst), .e(e), .q(q[4]) );
  my_DFF_1_3 fx_5 ( .d(d[5]), .clk(clk), .rst(rst), .e(e), .q(q[5]) );
  my_DFF_1_2 fx_6 ( .d(d[6]), .clk(clk), .rst(rst), .e(e), .q(q[6]) );
  my_DFF_1_1 fx_7 ( .d(d[7]), .clk(clk), .rst(rst), .e(e), .q(q[7]) );
endmodule


module reg_file_1 ( clk, rst, R, W, SP_EN, Rs1, Rs2, Rd, data_sp, data, S1, S2
 );
  input [1:0] Rs1;
  input [1:0] Rs2;
  input [1:0] Rd;
  input [7:0] data_sp;
  input [7:0] data;
  output [7:0] S1;
  output [7:0] S2;
  input clk, rst, R, W, SP_EN;
  wire   N75, N76, N77, N78, N90, N91, N92, N93, N94, N95, N96, N97, N98, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] R0;
  wire   [7:0] R1;
  wire   [7:0] R2;
  wire   [7:0] R3;
  wire   [7:0] R3_in;

  LATCHX1 \R3_in_reg[7]  ( .CLK(N90), .D(N98), .Q(R3_in[7]) );
  LATCHX1 \R3_in_reg[6]  ( .CLK(N90), .D(N97), .Q(R3_in[6]) );
  LATCHX1 \R3_in_reg[5]  ( .CLK(N90), .D(N96), .Q(R3_in[5]) );
  LATCHX1 \R3_in_reg[4]  ( .CLK(N90), .D(N95), .Q(R3_in[4]) );
  LATCHX1 \R3_in_reg[3]  ( .CLK(N90), .D(N94), .Q(R3_in[3]) );
  LATCHX1 \R3_in_reg[2]  ( .CLK(N90), .D(N93), .Q(R3_in[2]) );
  LATCHX1 \R3_in_reg[1]  ( .CLK(N90), .D(N92), .Q(R3_in[1]) );
  LATCHX1 \R3_in_reg[0]  ( .CLK(N90), .D(N91), .Q(R3_in[0]) );
  AO221X1 U21 ( .IN1(R3[7]), .IN2(n17), .IN3(R0[7]), .IN4(n2), .IN5(n18), .Q(
        S2[7]) );
  AO22X1 U22 ( .IN1(R2[7]), .IN2(n3), .IN3(R1[7]), .IN4(n5), .Q(n18) );
  AO221X1 U23 ( .IN1(R3[6]), .IN2(n17), .IN3(R0[6]), .IN4(n2), .IN5(n19), .Q(
        S2[6]) );
  AO22X1 U24 ( .IN1(R2[6]), .IN2(n3), .IN3(R1[6]), .IN4(n5), .Q(n19) );
  AO221X1 U25 ( .IN1(R3[5]), .IN2(n17), .IN3(R0[5]), .IN4(n2), .IN5(n20), .Q(
        S2[5]) );
  AO22X1 U26 ( .IN1(R2[5]), .IN2(n3), .IN3(R1[5]), .IN4(n5), .Q(n20) );
  AO221X1 U27 ( .IN1(R3[4]), .IN2(n17), .IN3(R0[4]), .IN4(n2), .IN5(n21), .Q(
        S2[4]) );
  AO22X1 U28 ( .IN1(R2[4]), .IN2(n3), .IN3(R1[4]), .IN4(n5), .Q(n21) );
  AO221X1 U29 ( .IN1(R3[3]), .IN2(n17), .IN3(R0[3]), .IN4(n2), .IN5(n22), .Q(
        S2[3]) );
  AO22X1 U30 ( .IN1(R2[3]), .IN2(n3), .IN3(R1[3]), .IN4(n5), .Q(n22) );
  AO221X1 U31 ( .IN1(R3[2]), .IN2(n17), .IN3(R0[2]), .IN4(n2), .IN5(n23), .Q(
        S2[2]) );
  AO22X1 U32 ( .IN1(R2[2]), .IN2(n3), .IN3(R1[2]), .IN4(n5), .Q(n23) );
  AO221X1 U33 ( .IN1(R3[1]), .IN2(n17), .IN3(R0[1]), .IN4(n2), .IN5(n24), .Q(
        S2[1]) );
  AO22X1 U34 ( .IN1(R2[1]), .IN2(n3), .IN3(R1[1]), .IN4(n5), .Q(n24) );
  AO221X1 U35 ( .IN1(R3[0]), .IN2(n17), .IN3(R0[0]), .IN4(n2), .IN5(n25), .Q(
        S2[0]) );
  AO22X1 U36 ( .IN1(R2[0]), .IN2(n3), .IN3(R1[0]), .IN4(n5), .Q(n25) );
  AND4X1 U37 ( .IN1(R), .IN2(n28), .IN3(n26), .IN4(n27), .Q(n17) );
  NAND3X0 U38 ( .IN1(R), .IN2(n4), .IN3(Rs2[1]), .QN(n27) );
  NAND3X0 U39 ( .IN1(R), .IN2(n6), .IN3(Rs2[0]), .QN(n26) );
  NAND3X0 U40 ( .IN1(n4), .IN2(n6), .IN3(R), .QN(n28) );
  AO221X1 U41 ( .IN1(n29), .IN2(R3[7]), .IN3(n7), .IN4(R0[7]), .IN5(n30), .Q(
        S1[7]) );
  AO22X1 U42 ( .IN1(n8), .IN2(R2[7]), .IN3(n10), .IN4(R1[7]), .Q(n30) );
  AO221X1 U43 ( .IN1(n29), .IN2(R3[6]), .IN3(n7), .IN4(R0[6]), .IN5(n31), .Q(
        S1[6]) );
  AO22X1 U44 ( .IN1(n8), .IN2(R2[6]), .IN3(n10), .IN4(R1[6]), .Q(n31) );
  AO221X1 U45 ( .IN1(n29), .IN2(R3[5]), .IN3(n7), .IN4(R0[5]), .IN5(n32), .Q(
        S1[5]) );
  AO22X1 U46 ( .IN1(n8), .IN2(R2[5]), .IN3(n10), .IN4(R1[5]), .Q(n32) );
  AO221X1 U47 ( .IN1(n29), .IN2(R3[4]), .IN3(n7), .IN4(R0[4]), .IN5(n33), .Q(
        S1[4]) );
  AO22X1 U48 ( .IN1(n8), .IN2(R2[4]), .IN3(n10), .IN4(R1[4]), .Q(n33) );
  AO221X1 U49 ( .IN1(n29), .IN2(R3[3]), .IN3(n7), .IN4(R0[3]), .IN5(n34), .Q(
        S1[3]) );
  AO22X1 U50 ( .IN1(n8), .IN2(R2[3]), .IN3(n10), .IN4(R1[3]), .Q(n34) );
  AO221X1 U51 ( .IN1(n29), .IN2(R3[2]), .IN3(n7), .IN4(R0[2]), .IN5(n35), .Q(
        S1[2]) );
  AO22X1 U52 ( .IN1(n8), .IN2(R2[2]), .IN3(n10), .IN4(R1[2]), .Q(n35) );
  AO221X1 U53 ( .IN1(n29), .IN2(R3[1]), .IN3(n7), .IN4(R0[1]), .IN5(n36), .Q(
        S1[1]) );
  AO22X1 U54 ( .IN1(n8), .IN2(R2[1]), .IN3(n10), .IN4(R1[1]), .Q(n36) );
  AO221X1 U55 ( .IN1(n29), .IN2(R3[0]), .IN3(n7), .IN4(R0[0]), .IN5(n37), .Q(
        S1[0]) );
  AO22X1 U56 ( .IN1(n8), .IN2(R2[0]), .IN3(n10), .IN4(R1[0]), .Q(n37) );
  AND4X1 U57 ( .IN1(R), .IN2(n40), .IN3(n38), .IN4(n39), .Q(n29) );
  NAND3X0 U58 ( .IN1(R), .IN2(n9), .IN3(Rs1[1]), .QN(n39) );
  NAND3X0 U59 ( .IN1(R), .IN2(n11), .IN3(Rs1[0]), .QN(n38) );
  NAND3X0 U60 ( .IN1(n9), .IN2(n11), .IN3(R), .QN(n40) );
  AO221X1 U61 ( .IN1(data_sp[7]), .IN2(n41), .IN3(data[7]), .IN4(n13), .IN5(
        rst), .Q(N98) );
  AO221X1 U62 ( .IN1(data_sp[6]), .IN2(n41), .IN3(data[6]), .IN4(n13), .IN5(
        rst), .Q(N97) );
  AO221X1 U63 ( .IN1(data_sp[5]), .IN2(n41), .IN3(data[5]), .IN4(n13), .IN5(
        rst), .Q(N96) );
  AO221X1 U64 ( .IN1(data_sp[4]), .IN2(n41), .IN3(data[4]), .IN4(n13), .IN5(
        rst), .Q(N95) );
  AO221X1 U65 ( .IN1(data_sp[3]), .IN2(n41), .IN3(data[3]), .IN4(n13), .IN5(
        rst), .Q(N94) );
  AO221X1 U66 ( .IN1(data_sp[2]), .IN2(n41), .IN3(data[2]), .IN4(n13), .IN5(
        rst), .Q(N93) );
  AO221X1 U67 ( .IN1(data_sp[1]), .IN2(n41), .IN3(data[1]), .IN4(n13), .IN5(
        rst), .Q(N92) );
  AO221X1 U68 ( .IN1(data_sp[0]), .IN2(n41), .IN3(data[0]), .IN4(n13), .IN5(
        rst), .Q(N91) );
  NAND3X0 U69 ( .IN1(n15), .IN2(n1), .IN3(n41), .QN(N90) );
  NAND3X0 U70 ( .IN1(n15), .IN2(n1), .IN3(n42), .QN(N78) );
  NAND3X0 U71 ( .IN1(Rd[1]), .IN2(Rd[0]), .IN3(W), .QN(n42) );
  NOR3X0 U72 ( .IN1(n43), .IN2(Rd[0]), .IN3(n14), .QN(N77) );
  NOR3X0 U73 ( .IN1(n43), .IN2(Rd[1]), .IN3(n12), .QN(N76) );
  NOR3X0 U74 ( .IN1(n43), .IN2(Rd[1]), .IN3(Rd[0]), .QN(N75) );
  my_nDFF_n8_4 R0_dest ( .clk(n16), .rst(rst), .e(N75), .d(data), .q(R0) );
  my_nDFF_n8_3 R1_dest ( .clk(n16), .rst(rst), .e(N76), .d(data), .q(R1) );
  my_nDFF_n8_2 R2_dest ( .clk(n16), .rst(rst), .e(N77), .d(data), .q(R2) );
  my_nDFF_n8_1 R3_dest ( .clk(n16), .rst(1'b0), .e(N78), .d(R3_in), .q(R3) );
  INVX0 U3 ( .IN(Rs1[1]), .QN(n11) );
  INVX0 U4 ( .IN(Rs1[0]), .QN(n9) );
  INVX0 U5 ( .IN(rst), .QN(n1) );
  NAND2X0 U6 ( .IN1(W), .IN2(n1), .QN(n43) );
  INVX0 U7 ( .IN(SP_EN), .QN(n15) );
  INVX0 U8 ( .IN(n40), .QN(n7) );
  INVX0 U9 ( .IN(n39), .QN(n8) );
  INVX0 U10 ( .IN(n38), .QN(n10) );
  INVX0 U11 ( .IN(n28), .QN(n2) );
  INVX0 U12 ( .IN(n26), .QN(n5) );
  INVX0 U13 ( .IN(n27), .QN(n3) );
  INVX0 U14 ( .IN(n41), .QN(n13) );
  INVX0 U15 ( .IN(Rd[1]), .QN(n14) );
  INVX0 U16 ( .IN(Rd[0]), .QN(n12) );
  INVX0 U17 ( .IN(Rs2[1]), .QN(n6) );
  INVX0 U18 ( .IN(Rs2[0]), .QN(n4) );
  NAND2X0 U19 ( .IN1(Rd[1]), .IN2(Rd[0]), .QN(n41) );
  INVX0 U20 ( .IN(clk), .QN(n16) );
endmodule


module my_DFF_1_164 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_163 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_162 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_161 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_160 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_159 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_158 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_157 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_156 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_155 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_154 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_153 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(d), .IN4(e), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_152 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4, n5, n6;

  DFFARX1 q_reg ( .D(n6), .CLK(clk), .RSTB(n5), .Q(q), .QN(n1) );
  INVX0 U2 ( .IN(rst), .QN(n5) );
  OR2X1 U3 ( .IN1(n1), .IN2(e), .Q(n2) );
  NAND2X0 U4 ( .IN1(e), .IN2(d), .QN(n4) );
  NAND2X0 U5 ( .IN1(n2), .IN2(n4), .QN(n6) );
endmodule


module my_DFF_1_151 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(d), .IN4(e), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_150 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_149 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_148 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_147 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_146 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_145 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_144 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_143 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_142 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_141 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_140 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_139 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_138 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_137 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_136 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_135 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_134 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_133 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_132 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_131 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_130 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_129 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_128 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_127 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_126 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_125 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_124 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_123 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_122 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_121 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_120 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_119 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_118 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_117 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_116 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_115 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_114 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_113 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_112 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_111 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_110 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_109 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_108 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_107 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_106 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_105 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_104 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_103 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_102 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_DFF_1_101 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n2), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n1), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n2) );
  INVX0 U4 ( .IN(e), .QN(n1) );
endmodule


module my_nDFF_n64 ( clk, rst, e, d, q );
  input [63:0] d;
  output [63:0] q;
  input clk, rst, e;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;

  my_DFF_1_164 fx_0 ( .d(d[0]), .clk(clk), .rst(n14), .e(n6), .q(q[0]) );
  my_DFF_1_163 fx_1 ( .d(d[1]), .clk(clk), .rst(n14), .e(n6), .q(q[1]) );
  my_DFF_1_162 fx_2 ( .d(d[2]), .clk(clk), .rst(n14), .e(n6), .q(q[2]) );
  my_DFF_1_161 fx_3 ( .d(d[3]), .clk(clk), .rst(n14), .e(n6), .q(q[3]) );
  my_DFF_1_160 fx_4 ( .d(d[4]), .clk(clk), .rst(n13), .e(n5), .q(q[4]) );
  my_DFF_1_159 fx_5 ( .d(d[5]), .clk(clk), .rst(n13), .e(n5), .q(q[5]) );
  my_DFF_1_158 fx_6 ( .d(d[6]), .clk(clk), .rst(n13), .e(n5), .q(q[6]) );
  my_DFF_1_157 fx_7 ( .d(d[7]), .clk(clk), .rst(n13), .e(n5), .q(q[7]) );
  my_DFF_1_156 fx_8 ( .d(d[8]), .clk(clk), .rst(n13), .e(n5), .q(q[8]) );
  my_DFF_1_155 fx_9 ( .d(d[9]), .clk(clk), .rst(n13), .e(n5), .q(q[9]) );
  my_DFF_1_154 fx_10 ( .d(d[10]), .clk(clk), .rst(n13), .e(n5), .q(q[10]) );
  my_DFF_1_153 fx_11 ( .d(d[11]), .clk(clk), .rst(n13), .e(n5), .q(q[11]) );
  my_DFF_1_152 fx_12 ( .d(d[12]), .clk(clk), .rst(n13), .e(n5), .q(q[12]) );
  my_DFF_1_151 fx_13 ( .d(d[13]), .clk(clk), .rst(n13), .e(n5), .q(q[13]) );
  my_DFF_1_150 fx_14 ( .d(d[14]), .clk(clk), .rst(n13), .e(n5), .q(q[14]) );
  my_DFF_1_149 fx_15 ( .d(d[15]), .clk(clk), .rst(n13), .e(n5), .q(q[15]) );
  my_DFF_1_148 fx_16 ( .d(d[16]), .clk(clk), .rst(n12), .e(n4), .q(q[16]) );
  my_DFF_1_147 fx_17 ( .d(d[17]), .clk(clk), .rst(n12), .e(n4), .q(q[17]) );
  my_DFF_1_146 fx_18 ( .d(d[18]), .clk(clk), .rst(n12), .e(n4), .q(q[18]) );
  my_DFF_1_145 fx_19 ( .d(d[19]), .clk(clk), .rst(n12), .e(n4), .q(q[19]) );
  my_DFF_1_144 fx_20 ( .d(d[20]), .clk(clk), .rst(n12), .e(n4), .q(q[20]) );
  my_DFF_1_143 fx_21 ( .d(d[21]), .clk(clk), .rst(n12), .e(n4), .q(q[21]) );
  my_DFF_1_142 fx_22 ( .d(d[22]), .clk(clk), .rst(n12), .e(n4), .q(q[22]) );
  my_DFF_1_141 fx_23 ( .d(d[23]), .clk(clk), .rst(n12), .e(n4), .q(q[23]) );
  my_DFF_1_140 fx_24 ( .d(d[24]), .clk(clk), .rst(n12), .e(n4), .q(q[24]) );
  my_DFF_1_139 fx_25 ( .d(d[25]), .clk(clk), .rst(n12), .e(n4), .q(q[25]) );
  my_DFF_1_138 fx_26 ( .d(d[26]), .clk(clk), .rst(n12), .e(n4), .q(q[26]) );
  my_DFF_1_137 fx_27 ( .d(d[27]), .clk(clk), .rst(n12), .e(n4), .q(q[27]) );
  my_DFF_1_136 fx_28 ( .d(d[28]), .clk(clk), .rst(n11), .e(n3), .q(q[28]) );
  my_DFF_1_135 fx_29 ( .d(d[29]), .clk(clk), .rst(n11), .e(n3), .q(q[29]) );
  my_DFF_1_134 fx_30 ( .d(d[30]), .clk(clk), .rst(n11), .e(n3), .q(q[30]) );
  my_DFF_1_133 fx_31 ( .d(d[31]), .clk(clk), .rst(n11), .e(n3), .q(q[31]) );
  my_DFF_1_132 fx_32 ( .d(d[32]), .clk(clk), .rst(n11), .e(n3), .q(q[32]) );
  my_DFF_1_131 fx_33 ( .d(d[33]), .clk(clk), .rst(n11), .e(n3), .q(q[33]) );
  my_DFF_1_130 fx_34 ( .d(d[34]), .clk(clk), .rst(n11), .e(n3), .q(q[34]) );
  my_DFF_1_129 fx_35 ( .d(d[35]), .clk(clk), .rst(n11), .e(n3), .q(q[35]) );
  my_DFF_1_128 fx_36 ( .d(d[36]), .clk(clk), .rst(n11), .e(n3), .q(q[36]) );
  my_DFF_1_127 fx_37 ( .d(d[37]), .clk(clk), .rst(n11), .e(n3), .q(q[37]) );
  my_DFF_1_126 fx_38 ( .d(d[38]), .clk(clk), .rst(n11), .e(n3), .q(q[38]) );
  my_DFF_1_125 fx_39 ( .d(d[39]), .clk(clk), .rst(n11), .e(n3), .q(q[39]) );
  my_DFF_1_124 fx_40 ( .d(d[40]), .clk(clk), .rst(n10), .e(n2), .q(q[40]) );
  my_DFF_1_123 fx_41 ( .d(d[41]), .clk(clk), .rst(n10), .e(n2), .q(q[41]) );
  my_DFF_1_122 fx_42 ( .d(d[42]), .clk(clk), .rst(n10), .e(n2), .q(q[42]) );
  my_DFF_1_121 fx_43 ( .d(d[43]), .clk(clk), .rst(n10), .e(n2), .q(q[43]) );
  my_DFF_1_120 fx_44 ( .d(d[44]), .clk(clk), .rst(n10), .e(n2), .q(q[44]) );
  my_DFF_1_119 fx_45 ( .d(d[45]), .clk(clk), .rst(n10), .e(n2), .q(q[45]) );
  my_DFF_1_118 fx_46 ( .d(d[46]), .clk(clk), .rst(n10), .e(n2), .q(q[46]) );
  my_DFF_1_117 fx_47 ( .d(d[47]), .clk(clk), .rst(n10), .e(n2), .q(q[47]) );
  my_DFF_1_116 fx_48 ( .d(d[48]), .clk(clk), .rst(n10), .e(n2), .q(q[48]) );
  my_DFF_1_115 fx_49 ( .d(d[49]), .clk(clk), .rst(n10), .e(n2), .q(q[49]) );
  my_DFF_1_114 fx_50 ( .d(d[50]), .clk(clk), .rst(n10), .e(n2), .q(q[50]) );
  my_DFF_1_113 fx_51 ( .d(d[51]), .clk(clk), .rst(n10), .e(n2), .q(q[51]) );
  my_DFF_1_112 fx_52 ( .d(d[52]), .clk(clk), .rst(n9), .e(n1), .q(q[52]) );
  my_DFF_1_111 fx_53 ( .d(d[53]), .clk(clk), .rst(n9), .e(n1), .q(q[53]) );
  my_DFF_1_110 fx_54 ( .d(d[54]), .clk(clk), .rst(n9), .e(n1), .q(q[54]) );
  my_DFF_1_109 fx_55 ( .d(d[55]), .clk(clk), .rst(n9), .e(n1), .q(q[55]) );
  my_DFF_1_108 fx_56 ( .d(d[56]), .clk(clk), .rst(n9), .e(n1), .q(q[56]) );
  my_DFF_1_107 fx_57 ( .d(d[57]), .clk(clk), .rst(n9), .e(n1), .q(q[57]) );
  my_DFF_1_106 fx_58 ( .d(d[58]), .clk(clk), .rst(n9), .e(n1), .q(q[58]) );
  my_DFF_1_105 fx_59 ( .d(d[59]), .clk(clk), .rst(n9), .e(n1), .q(q[59]) );
  my_DFF_1_104 fx_60 ( .d(d[60]), .clk(clk), .rst(n9), .e(n1), .q(q[60]) );
  my_DFF_1_103 fx_61 ( .d(d[61]), .clk(clk), .rst(n9), .e(n1), .q(q[61]) );
  my_DFF_1_102 fx_62 ( .d(d[62]), .clk(clk), .rst(n9), .e(n1), .q(q[62]) );
  my_DFF_1_101 fx_63 ( .d(d[63]), .clk(clk), .rst(n9), .e(n1), .q(q[63]) );
  NBUFFX2 U1 ( .IN(n7), .Q(n5) );
  NBUFFX2 U2 ( .IN(n7), .Q(n4) );
  NBUFFX2 U3 ( .IN(n8), .Q(n3) );
  NBUFFX2 U4 ( .IN(n8), .Q(n2) );
  NBUFFX2 U5 ( .IN(n8), .Q(n1) );
  NBUFFX2 U6 ( .IN(n7), .Q(n6) );
  NBUFFX2 U7 ( .IN(n15), .Q(n13) );
  NBUFFX2 U8 ( .IN(n15), .Q(n12) );
  NBUFFX2 U9 ( .IN(n16), .Q(n11) );
  NBUFFX2 U10 ( .IN(n16), .Q(n10) );
  NBUFFX2 U11 ( .IN(n16), .Q(n9) );
  NBUFFX2 U12 ( .IN(n15), .Q(n14) );
  NBUFFX2 U13 ( .IN(e), .Q(n7) );
  NBUFFX2 U14 ( .IN(e), .Q(n8) );
  NBUFFX2 U15 ( .IN(rst), .Q(n15) );
  NBUFFX2 U16 ( .IN(rst), .Q(n16) );
endmodule


module my_adder_1_0 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n1, n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(n1), .IN4(cin), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n1) );
  NBUFFX2 U4 ( .IN(n1), .Q(n2) );
endmodule


module my_adder_1_15 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_14 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2, n3;

  XOR2X1 U1 ( .IN1(n2), .IN2(n3), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n3), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n3) );
  NBUFFX2 U4 ( .IN(cin), .Q(n2) );
endmodule


module my_adder_1_13 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2, n3;

  XOR2X1 U1 ( .IN1(n2), .IN2(n3), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n3), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n3) );
  NBUFFX2 U4 ( .IN(cin), .Q(n2) );
endmodule


module my_adder_1_12 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_11 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2, n3, n4;

  XOR2X1 U1 ( .IN1(n3), .IN2(n4), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n4), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n4) );
  INVX0 U4 ( .IN(cin), .QN(n2) );
  INVX0 U5 ( .IN(n2), .QN(n3) );
endmodule


module my_adder_1_10 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_9 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(n2), .IN2(cin), .Q(s) );
  XOR2X1 U3 ( .IN1(b), .IN2(a), .Q(n2) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
endmodule


module my_nadder_n8_0 ( a, b, cin, s, cout );
  input [7:0] a;
  input [7:0] b;
  output [7:0] s;
  input cin;
  output cout;

  wire   [6:0] temp;

  my_adder_1_0 f0 ( .a(a[0]), .b(b[0]), .cin(cin), .s(s[0]), .cout(temp[0]) );
  my_adder_1_15 fx_1 ( .a(a[1]), .b(b[1]), .cin(temp[0]), .s(s[1]), .cout(
        temp[1]) );
  my_adder_1_14 fx_2 ( .a(a[2]), .b(b[2]), .cin(temp[1]), .s(s[2]), .cout(
        temp[2]) );
  my_adder_1_13 fx_3 ( .a(a[3]), .b(b[3]), .cin(temp[2]), .s(s[3]), .cout(
        temp[3]) );
  my_adder_1_12 fx_4 ( .a(a[4]), .b(b[4]), .cin(temp[3]), .s(s[4]), .cout(
        temp[4]) );
  my_adder_1_11 fx_5 ( .a(a[5]), .b(b[5]), .cin(temp[4]), .s(s[5]), .cout(
        temp[5]) );
  my_adder_1_10 fx_6 ( .a(a[6]), .b(b[6]), .cin(temp[5]), .s(s[6]), .cout(
        temp[6]) );
  my_adder_1_9 fx_7 ( .a(a[7]), .b(b[7]), .cin(temp[6]), .s(s[7]), .cout(cout)
         );
endmodule


module partA_1 ( a, b, s, F, cout, zero, negative, overflow );
  input [7:0] a;
  input [7:0] b;
  output [7:0] F;
  input s;
  output cout, zero, negative, overflow;
  wire   n10, N17, N18, N19, N20, N21, N22, N23, N24, cout1, N25, n4, n5, n6,
         n7, n1, n3, n8, n9;
  assign negative = F[7];
  assign overflow = N25;

  OR4X1 U6 ( .IN1(F[1]), .IN2(F[0]), .IN3(F[3]), .IN4(F[2]), .Q(n5) );
  OR4X1 U7 ( .IN1(F[5]), .IN2(F[4]), .IN3(n10), .IN4(F[6]), .Q(n4) );
  XNOR2X1 U8 ( .IN1(n3), .IN2(cout1), .Q(cout) );
  XOR2X1 U11 ( .IN1(s), .IN2(b[7]), .Q(N24) );
  XNOR2X1 U12 ( .IN1(n3), .IN2(b[6]), .Q(N23) );
  XNOR2X1 U13 ( .IN1(n3), .IN2(b[5]), .Q(N22) );
  XNOR2X1 U14 ( .IN1(n3), .IN2(b[4]), .Q(N21) );
  XNOR2X1 U15 ( .IN1(n3), .IN2(b[3]), .Q(N20) );
  XNOR2X1 U16 ( .IN1(n3), .IN2(b[2]), .Q(N19) );
  XNOR2X1 U17 ( .IN1(n3), .IN2(b[1]), .Q(N18) );
  my_nadder_n8_0 u0 ( .a(a), .b({N24, N23, N22, N21, N20, N19, N18, N17}), 
        .cin(s), .s({n10, F[6:0]}), .cout(cout1) );
  INVX0 U1 ( .IN(n10), .QN(n1) );
  XOR2X1 U2 ( .IN1(s), .IN2(b[0]), .Q(N17) );
  INVX0 U3 ( .IN(n1), .QN(F[7]) );
  INVX0 U4 ( .IN(s), .QN(n3) );
  OR3X1 U5 ( .IN1(n9), .IN2(F[7]), .IN3(n8), .Q(n6) );
  NAND3X0 U9 ( .IN1(n9), .IN2(n8), .IN3(F[7]), .QN(n7) );
  INVX0 U10 ( .IN(a[7]), .QN(n8) );
  INVX0 U18 ( .IN(N24), .QN(n9) );
  NAND2X0 U19 ( .IN1(n6), .IN2(n7), .QN(N25) );
  NOR2X0 U20 ( .IN1(n4), .IN2(n5), .QN(zero) );
endmodule


module partB_1 ( a, b, s, F, zero, negative );
  input [7:0] a;
  input [7:0] b;
  output [7:0] F;
  input s;
  output zero, negative;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  assign F[0] = N18;
  assign F[1] = N19;
  assign F[2] = N20;
  assign F[3] = N21;
  assign F[4] = N22;
  assign F[5] = N23;
  assign F[6] = N24;
  assign negative = N25;
  assign F[7] = N25;

  OR4X1 U2 ( .IN1(N18), .IN2(N19), .IN3(N20), .IN4(N21), .Q(n2) );
  OR4X1 U3 ( .IN1(N22), .IN2(N23), .IN3(N24), .IN4(N25), .Q(n1) );
  AO22X1 U4 ( .IN1(b[7]), .IN2(a[7]), .IN3(n11), .IN4(n3), .Q(N25) );
  OR2X1 U5 ( .IN1(b[7]), .IN2(a[7]), .Q(n3) );
  AO22X1 U6 ( .IN1(b[6]), .IN2(a[6]), .IN3(n11), .IN4(n4), .Q(N24) );
  OR2X1 U7 ( .IN1(b[6]), .IN2(a[6]), .Q(n4) );
  AO22X1 U8 ( .IN1(b[5]), .IN2(a[5]), .IN3(n11), .IN4(n5), .Q(N23) );
  OR2X1 U9 ( .IN1(b[5]), .IN2(a[5]), .Q(n5) );
  AO22X1 U10 ( .IN1(b[4]), .IN2(a[4]), .IN3(n11), .IN4(n6), .Q(N22) );
  OR2X1 U11 ( .IN1(b[4]), .IN2(a[4]), .Q(n6) );
  AO22X1 U12 ( .IN1(b[3]), .IN2(a[3]), .IN3(n11), .IN4(n7), .Q(N21) );
  OR2X1 U13 ( .IN1(b[3]), .IN2(a[3]), .Q(n7) );
  AO22X1 U14 ( .IN1(b[2]), .IN2(a[2]), .IN3(n11), .IN4(n8), .Q(N20) );
  OR2X1 U15 ( .IN1(b[2]), .IN2(a[2]), .Q(n8) );
  AO22X1 U16 ( .IN1(b[1]), .IN2(a[1]), .IN3(n11), .IN4(n9), .Q(N19) );
  OR2X1 U17 ( .IN1(b[1]), .IN2(a[1]), .Q(n9) );
  AO22X1 U18 ( .IN1(b[0]), .IN2(a[0]), .IN3(n11), .IN4(n10), .Q(N18) );
  OR2X1 U19 ( .IN1(b[0]), .IN2(a[0]), .Q(n10) );
  NBUFFX2 U1 ( .IN(s), .Q(n11) );
  NOR2X0 U20 ( .IN1(n1), .IN2(n2), .QN(zero) );
endmodule


module partC_1 ( a, s, cin, F, Cout, zero, negative );
  input [7:0] a;
  output [7:0] F;
  input s, cin;
  output Cout, zero, negative;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, n2, n3, n4, n1, n5;
  assign F[0] = N2;
  assign F[1] = N3;
  assign F[2] = N4;
  assign F[3] = N5;
  assign F[4] = N6;
  assign F[5] = N7;
  assign F[6] = N8;
  assign negative = N9;
  assign F[7] = N9;
  assign Cout = N10;

  OA22X1 U3 ( .IN1(n1), .IN2(a[0]), .IN3(a[7]), .IN4(n5), .Q(n4) );
  OR2X1 U4 ( .IN1(a[2]), .IN2(a[3]), .Q(n3) );
  AO22X1 U6 ( .IN1(cin), .IN2(n1), .IN3(a[6]), .IN4(n5), .Q(N9) );
  AO22X1 U7 ( .IN1(a[7]), .IN2(n1), .IN3(a[5]), .IN4(n5), .Q(N8) );
  AO22X1 U8 ( .IN1(a[6]), .IN2(n1), .IN3(a[4]), .IN4(n5), .Q(N7) );
  AO22X1 U9 ( .IN1(a[5]), .IN2(n1), .IN3(a[3]), .IN4(n5), .Q(N6) );
  AO22X1 U10 ( .IN1(a[4]), .IN2(n1), .IN3(a[2]), .IN4(n5), .Q(N5) );
  AO22X1 U11 ( .IN1(a[3]), .IN2(n1), .IN3(a[1]), .IN4(n5), .Q(N4) );
  AO22X1 U12 ( .IN1(a[2]), .IN2(n1), .IN3(a[0]), .IN4(n5), .Q(N3) );
  AO22X1 U13 ( .IN1(cin), .IN2(n5), .IN3(a[1]), .IN4(n1), .Q(N2) );
  AO22X1 U14 ( .IN1(a[7]), .IN2(n5), .IN3(a[0]), .IN4(n1), .Q(N10) );
  INVX0 U1 ( .IN(n1), .QN(n5) );
  NBUFFX2 U2 ( .IN(s), .Q(n1) );
  OR4X1 U5 ( .IN1(a[4]), .IN2(a[5]), .IN3(a[6]), .IN4(cin), .Q(n2) );
  NOR4X0 U15 ( .IN1(n2), .IN2(n3), .IN3(a[1]), .IN4(n4), .QN(zero) );
endmodule


module my_adder_1_8 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(n2), .IN4(cin), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_7 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_6 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_5 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_4 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_3 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_2 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_adder_1_1 ( a, b, cin, s, cout );
  input a, b, cin;
  output s, cout;
  wire   n2;

  XOR2X1 U1 ( .IN1(cin), .IN2(n2), .Q(s) );
  AO22X1 U2 ( .IN1(a), .IN2(b), .IN3(cin), .IN4(n2), .Q(cout) );
  XOR2X1 U3 ( .IN1(a), .IN2(b), .Q(n2) );
endmodule


module my_nadder_n8_1 ( a, b, cin, s, cout );
  input [7:0] a;
  input [7:0] b;
  output [7:0] s;
  input cin;
  output cout;

  wire   [6:0] temp;

  my_adder_1_8 f0 ( .a(a[0]), .b(b[0]), .cin(cin), .s(s[0]), .cout(temp[0]) );
  my_adder_1_7 fx_1 ( .a(a[1]), .b(b[1]), .cin(temp[0]), .s(s[1]), .cout(
        temp[1]) );
  my_adder_1_6 fx_2 ( .a(a[2]), .b(b[2]), .cin(temp[1]), .s(s[2]), .cout(
        temp[2]) );
  my_adder_1_5 fx_3 ( .a(a[3]), .b(b[3]), .cin(temp[2]), .s(s[3]), .cout(
        temp[3]) );
  my_adder_1_4 fx_4 ( .a(a[4]), .b(b[4]), .cin(temp[3]), .s(s[4]), .cout(
        temp[4]) );
  my_adder_1_3 fx_5 ( .a(a[5]), .b(b[5]), .cin(temp[4]), .s(s[5]), .cout(
        temp[5]) );
  my_adder_1_2 fx_6 ( .a(a[6]), .b(b[6]), .cin(temp[5]), .s(s[6]), .cout(
        temp[6]) );
  my_adder_1_1 fx_7 ( .a(a[7]), .b(b[7]), .cin(temp[6]), .s(s[7]), .cout(cout)
         );
endmodule


module partD_1 ( a, s, F, Cout, zero, negative, overflow );
  input [7:0] a;
  input [1:0] s;
  output [7:0] F;
  output Cout, zero, negative, overflow;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, cin, cout_tmp, n5, n6, n7, n8,
         n9, n1, n2, n3, n4, n10;
  assign negative = F[7];

  OA22X1 U9 ( .IN1(n5), .IN2(n6), .IN3(a[7]), .IN4(n2), .Q(overflow) );
  AND3X1 U10 ( .IN1(n1), .IN2(n3), .IN3(F[7]), .Q(n5) );
  OR4X1 U11 ( .IN1(F[1]), .IN2(F[0]), .IN3(F[3]), .IN4(F[2]), .Q(n9) );
  OR4X1 U12 ( .IN1(F[7]), .IN2(F[4]), .IN3(F[5]), .IN4(F[6]), .Q(n8) );
  XNOR2X1 U13 ( .IN1(n10), .IN2(s[0]), .Q(cin) );
  XNOR2X1 U15 ( .IN1(n1), .IN2(a[6]), .Q(N17) );
  XNOR2X1 U16 ( .IN1(n1), .IN2(a[5]), .Q(N16) );
  XNOR2X1 U17 ( .IN1(n1), .IN2(a[4]), .Q(N15) );
  XNOR2X1 U18 ( .IN1(n1), .IN2(a[3]), .Q(N14) );
  XNOR2X1 U19 ( .IN1(n1), .IN2(a[2]), .Q(N13) );
  XNOR2X1 U20 ( .IN1(n1), .IN2(a[1]), .Q(N12) );
  XNOR2X1 U22 ( .IN1(cout_tmp), .IN2(n7), .Q(Cout) );
  my_nadder_n8_1 u0 ( .a({N18, N17, N16, N15, N14, N13, N12, N11}), .b({n4, n4, 
        n4, n4, n4, n4, n4, n4}), .cin(cin), .s(F), .cout(cout_tmp) );
  XOR2X1 U2 ( .IN1(a[0]), .IN2(n10), .Q(N11) );
  INVX0 U3 ( .IN(s[0]), .QN(n2) );
  INVX0 U4 ( .IN(n7), .QN(n4) );
  INVX0 U5 ( .IN(a[7]), .QN(n3) );
  NAND2X0 U6 ( .IN1(s[0]), .IN2(s[1]), .QN(n7) );
  NBUFFX2 U7 ( .IN(s[1]), .Q(n1) );
  XOR2X1 U8 ( .IN1(a[7]), .IN2(n10), .Q(N18) );
  INVX0 U14 ( .IN(n1), .QN(n10) );
  NOR2X0 U21 ( .IN1(F[7]), .IN2(n7), .QN(n6) );
  NOR2X0 U23 ( .IN1(n8), .IN2(n9), .QN(zero) );
endmodule


module ALSU ( a, b, s, cin, F, cout, zero, negative, overflow );
  input [7:0] a;
  input [7:0] b;
  input [3:0] s;
  output [7:0] F;
  input cin;
  output cout, zero, negative, overflow;
  wire   N57, N58, N59, N60, N61, N62, N63, N64, N65, n1, n2, n3, n4, n5, n8,
         n10, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n6, n7, n9, n11, n12, n32;
  wire   [7:0] w0;
  wire   [2:0] carries;
  wire   [3:0] zeros;
  wire   [3:0] negatives;
  wire   [1:0] overflows;
  wire   [7:0] w1;
  wire   [7:0] w2;
  wire   [7:0] w3;
  tri   cout;
  tri   zero;
  tri   negative;
  tri   overflow;

  LATCHX1 \F_reg[7]  ( .CLK(N57), .D(N65), .Q(F[7]) );
  LATCHX1 \F_reg[6]  ( .CLK(N57), .D(N64), .Q(F[6]) );
  LATCHX1 \F_reg[5]  ( .CLK(N57), .D(N63), .Q(F[5]) );
  LATCHX1 \F_reg[4]  ( .CLK(N57), .D(N62), .Q(F[4]) );
  LATCHX1 \F_reg[3]  ( .CLK(N57), .D(N61), .Q(F[3]) );
  LATCHX1 \F_reg[2]  ( .CLK(N57), .D(N60), .Q(F[2]) );
  LATCHX1 \F_reg[1]  ( .CLK(N57), .D(N59), .Q(F[1]) );
  LATCHX1 \F_reg[0]  ( .CLK(N57), .D(N58), .Q(F[0]) );
  TNBUFFX1 overflow_tri ( .INP(n31), .ENB(n29), .Z(overflow) );
  TNBUFFX1 negative_tri ( .INP(n30), .ENB(n29), .Z(negative) );
  TNBUFFX1 cout_tri ( .INP(n26), .ENB(n27), .Z(cout) );
  AO221X1 U3 ( .IN1(zeros[1]), .IN2(n1), .IN3(zeros[2]), .IN4(n2), .IN5(n3), 
        .Q(n28) );
  AO22X1 U4 ( .IN1(zeros[3]), .IN2(s[3]), .IN3(zeros[0]), .IN4(n4), .Q(n3) );
  AO22X1 U5 ( .IN1(overflows[1]), .IN2(s[3]), .IN3(overflows[0]), .IN4(n4), 
        .Q(n31) );
  AO221X1 U6 ( .IN1(negatives[1]), .IN2(n1), .IN3(negatives[2]), .IN4(n2), 
        .IN5(n5), .Q(n30) );
  AO22X1 U7 ( .IN1(negatives[3]), .IN2(s[3]), .IN3(negatives[0]), .IN4(n4), 
        .Q(n5) );
  AOI21X1 U8 ( .IN1(n4), .IN2(n9), .IN3(n12), .QN(n29) );
  AO221X1 U9 ( .IN1(carries[2]), .IN2(n8), .IN3(n12), .IN4(n7), .IN5(n10), .Q(
        n26) );
  AO22X1 U10 ( .IN1(carries[0]), .IN2(n4), .IN3(carries[1]), .IN4(n2), .Q(n10)
         );
  AO222X1 U13 ( .IN1(s[1]), .IN2(n11), .IN3(s[3]), .IN4(n9), .IN5(s[2]), .IN6(
        n32), .Q(n27) );
  AO222X1 U15 ( .IN1(w1[7]), .IN2(n16), .IN3(w2[7]), .IN4(n17), .IN5(w3[7]), 
        .IN6(n8), .Q(n15) );
  AO222X1 U17 ( .IN1(w1[6]), .IN2(n16), .IN3(w2[6]), .IN4(n17), .IN5(w3[6]), 
        .IN6(n8), .Q(n18) );
  AO221X1 U18 ( .IN1(w0[5]), .IN2(n13), .IN3(b[5]), .IN4(n14), .IN5(n19), .Q(
        N63) );
  AO222X1 U19 ( .IN1(w1[5]), .IN2(n16), .IN3(w2[5]), .IN4(n17), .IN5(w3[5]), 
        .IN6(n8), .Q(n19) );
  AO221X1 U20 ( .IN1(w0[4]), .IN2(n13), .IN3(b[4]), .IN4(n14), .IN5(n20), .Q(
        N62) );
  AO222X1 U21 ( .IN1(w1[4]), .IN2(n16), .IN3(w2[4]), .IN4(n17), .IN5(w3[4]), 
        .IN6(n8), .Q(n20) );
  AO221X1 U22 ( .IN1(w0[3]), .IN2(n13), .IN3(b[3]), .IN4(n14), .IN5(n21), .Q(
        N61) );
  AO222X1 U23 ( .IN1(w1[3]), .IN2(n16), .IN3(w2[3]), .IN4(n17), .IN5(w3[3]), 
        .IN6(n8), .Q(n21) );
  AO221X1 U24 ( .IN1(w0[2]), .IN2(n13), .IN3(b[2]), .IN4(n14), .IN5(n22), .Q(
        N60) );
  AO222X1 U25 ( .IN1(w1[2]), .IN2(n16), .IN3(w2[2]), .IN4(n17), .IN5(w3[2]), 
        .IN6(n8), .Q(n22) );
  AO221X1 U26 ( .IN1(w0[1]), .IN2(n13), .IN3(b[1]), .IN4(n14), .IN5(n23), .Q(
        N59) );
  AO222X1 U27 ( .IN1(w1[1]), .IN2(n16), .IN3(w2[1]), .IN4(n17), .IN5(w3[1]), 
        .IN6(n8), .Q(n23) );
  AO221X1 U28 ( .IN1(w0[0]), .IN2(n13), .IN3(n6), .IN4(n14), .IN5(n24), .Q(N58) );
  AO222X1 U29 ( .IN1(w1[0]), .IN2(n16), .IN3(w2[0]), .IN4(n17), .IN5(w3[0]), 
        .IN6(n8), .Q(n24) );
  AND2X1 U31 ( .IN1(n2), .IN2(n32), .Q(n17) );
  AND2X1 U35 ( .IN1(s[2]), .IN2(n1), .Q(n16) );
  NAND3X0 U38 ( .IN1(n4), .IN2(n9), .IN3(s[0]), .QN(n25) );
  AND2X1 U40 ( .IN1(n4), .IN2(s[1]), .Q(n13) );
  partA_1 u0 ( .a(a), .b(b), .s(s[0]), .F(w0), .cout(carries[0]), .zero(
        zeros[0]), .negative(negatives[0]), .overflow(overflows[0]) );
  partB_1 u1 ( .a(a), .b({b[7:1], n6}), .s(s[0]), .F(w1), .zero(zeros[1]), 
        .negative(negatives[1]) );
  partC_1 u2 ( .a({b[7:1], n6}), .s(s[0]), .cin(cin), .F(w2), .Cout(carries[1]), .zero(zeros[2]), .negative(negatives[2]) );
  partD_1 u3 ( .a(b), .s(s[1:0]), .F(w3), .Cout(carries[2]), .zero(zeros[3]), 
        .negative(negatives[3]), .overflow(overflows[1]) );
  TNBUFFX2 zero_tri ( .INP(n28), .ENB(n29), .Z(zero) );
  NBUFFX2 U11 ( .IN(b[0]), .Q(n6) );
  NOR2X0 U12 ( .IN1(n11), .IN2(n9), .QN(n2) );
  INVX0 U14 ( .IN(N57), .QN(n12) );
  AO221X1 U16 ( .IN1(w0[6]), .IN2(n13), .IN3(b[6]), .IN4(n14), .IN5(n18), .Q(
        N64) );
  AO221X1 U30 ( .IN1(w0[7]), .IN2(n13), .IN3(b[7]), .IN4(n14), .IN5(n15), .Q(
        N65) );
  NAND2X0 U32 ( .IN1(N57), .IN2(n25), .QN(n14) );
  INVX0 U33 ( .IN(s[0]), .QN(n7) );
  NOR2X0 U34 ( .IN1(s[2]), .IN2(s[3]), .QN(n4) );
  NAND2X0 U36 ( .IN1(s[3]), .IN2(s[2]), .QN(N57) );
  INVX0 U37 ( .IN(s[1]), .QN(n9) );
  NOR2X0 U39 ( .IN1(s[1]), .IN2(s[3]), .QN(n1) );
  INVX0 U41 ( .IN(s[2]), .QN(n11) );
  NOR2X0 U42 ( .IN1(n32), .IN2(s[2]), .QN(n8) );
  INVX0 U43 ( .IN(s[3]), .QN(n32) );
endmodule


module execute_1 ( ID_EX, flags_in, mem_data, mem_rd, mem_acc_mode, stall_Rd, 
        mem_valid, wb_data, wb_rd, wb_valid, sp_data, sp_en, IN_PORT, EX_MEM, 
        flags_out, stall, ret_ex, branch, target_addr, rti );
  input [63:0] ID_EX;
  input [3:0] flags_in;
  input [7:0] mem_data;
  input [1:0] mem_rd;
  input [2:0] mem_acc_mode;
  input [1:0] stall_Rd;
  input [7:0] wb_data;
  input [1:0] wb_rd;
  input [7:0] sp_data;
  input [7:0] IN_PORT;
  output [31:0] EX_MEM;
  output [3:0] flags_out;
  output [7:0] target_addr;
  input mem_valid, wb_valid, sp_en;
  output stall, ret_ex, branch, rti;
  wire   ID_EX_56, ID_EX_55, ID_EX_54, ID_EX_53, ID_EX_52, ID_EX_51, ID_EX_50,
         ID_EX_49, ID_EX_48, ID_EX_47, ID_EX_46, ID_EX_45, ID_EX_44, ID_EX_43,
         ID_EX_41, ID_EX_40, ID_EX_39, ID_EX_38, ID_EX_34, \ID_EX[57] ,
         \ID_EX[42] , \ID_EX[37] , \ID_EX[36] , \ID_EX[35] , \ID_EX[33] ,
         \ID_EX[32] , N120, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n119,
         n120, n121, n122, n123, n124, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31;
  wire   [7:0] s1_tmp;
  wire   [7:0] alu_b;
  wire   [7:0] result;
  tri   [3:0] CCR;
  assign EX_MEM[24] = 1'b0;
  assign EX_MEM[25] = 1'b0;
  assign EX_MEM[26] = 1'b0;
  assign EX_MEM[27] = 1'b0;
  assign EX_MEM[28] = 1'b0;
  assign EX_MEM[29] = 1'b0;
  assign EX_MEM[30] = 1'b0;
  assign EX_MEM[31] = 1'b0;
  assign rti = ID_EX_56;
  assign ID_EX_56 = ID_EX[56];
  assign ID_EX_55 = ID_EX[55];
  assign ID_EX_54 = ID_EX[54];
  assign ID_EX_53 = ID_EX[53];
  assign ID_EX_52 = ID_EX[52];
  assign ID_EX_51 = ID_EX[51];
  assign ID_EX_50 = ID_EX[50];
  assign ID_EX_49 = ID_EX[49];
  assign ID_EX_48 = ID_EX[48];
  assign ID_EX_47 = ID_EX[47];
  assign ID_EX_46 = ID_EX[46];
  assign ID_EX_45 = ID_EX[45];
  assign ID_EX_44 = ID_EX[44];
  assign ID_EX_43 = ID_EX[43];
  assign ID_EX_41 = ID_EX[41];
  assign ID_EX_40 = ID_EX[40];
  assign ID_EX_39 = ID_EX[39];
  assign ID_EX_38 = ID_EX[38];
  assign ID_EX_34 = ID_EX[34];
  assign EX_MEM[23] = \ID_EX[57] ;
  assign \ID_EX[57]  = ID_EX[57];
  assign ret_ex = \ID_EX[42] ;
  assign EX_MEM[22] = \ID_EX[42] ;
  assign \ID_EX[42]  = ID_EX[42];
  assign EX_MEM[20] = \ID_EX[37] ;
  assign \ID_EX[37]  = ID_EX[37];
  assign EX_MEM[19] = \ID_EX[36] ;
  assign \ID_EX[36]  = ID_EX[36];
  assign EX_MEM[18] = \ID_EX[35] ;
  assign \ID_EX[35]  = ID_EX[35];
  assign EX_MEM[17] = \ID_EX[33] ;
  assign \ID_EX[33]  = ID_EX[33];
  assign EX_MEM[16] = \ID_EX[32] ;
  assign \ID_EX[32]  = ID_EX[32];
  assign stall = N120;

  AO221X1 U43 ( .IN1(ID_EX_55), .IN2(n44), .IN3(sp_data[7]), .IN4(n45), .IN5(
        n46), .Q(target_addr[7]) );
  AO22X1 U44 ( .IN1(mem_data[7]), .IN2(n47), .IN3(wb_data[7]), .IN4(n48), .Q(
        n46) );
  AO221X1 U45 ( .IN1(ID_EX_54), .IN2(n44), .IN3(sp_data[6]), .IN4(n45), .IN5(
        n49), .Q(target_addr[6]) );
  AO22X1 U46 ( .IN1(mem_data[6]), .IN2(n47), .IN3(wb_data[6]), .IN4(n48), .Q(
        n49) );
  AO221X1 U47 ( .IN1(ID_EX_53), .IN2(n44), .IN3(sp_data[5]), .IN4(n45), .IN5(
        n50), .Q(target_addr[5]) );
  AO22X1 U48 ( .IN1(mem_data[5]), .IN2(n47), .IN3(wb_data[5]), .IN4(n48), .Q(
        n50) );
  AO221X1 U49 ( .IN1(ID_EX_52), .IN2(n44), .IN3(sp_data[4]), .IN4(n45), .IN5(
        n51), .Q(target_addr[4]) );
  AO22X1 U50 ( .IN1(mem_data[4]), .IN2(n47), .IN3(wb_data[4]), .IN4(n48), .Q(
        n51) );
  AO221X1 U51 ( .IN1(ID_EX_51), .IN2(n44), .IN3(sp_data[3]), .IN4(n45), .IN5(
        n52), .Q(target_addr[3]) );
  AO22X1 U52 ( .IN1(mem_data[3]), .IN2(n47), .IN3(wb_data[3]), .IN4(n48), .Q(
        n52) );
  AO221X1 U53 ( .IN1(ID_EX_50), .IN2(n44), .IN3(sp_data[2]), .IN4(n45), .IN5(
        n53), .Q(target_addr[2]) );
  AO22X1 U54 ( .IN1(mem_data[2]), .IN2(n47), .IN3(wb_data[2]), .IN4(n48), .Q(
        n53) );
  AO221X1 U55 ( .IN1(ID_EX_49), .IN2(n44), .IN3(sp_data[1]), .IN4(n45), .IN5(
        n54), .Q(target_addr[1]) );
  AO22X1 U56 ( .IN1(mem_data[1]), .IN2(n47), .IN3(wb_data[1]), .IN4(n48), .Q(
        n54) );
  AO221X1 U57 ( .IN1(ID_EX_48), .IN2(n44), .IN3(sp_data[0]), .IN4(n45), .IN5(
        n55), .Q(target_addr[0]) );
  AO22X1 U58 ( .IN1(mem_data[0]), .IN2(n47), .IN3(wb_data[0]), .IN4(n48), .Q(
        n55) );
  AND2X1 U59 ( .IN1(n57), .IN2(n56), .Q(n44) );
  NAND3X0 U60 ( .IN1(ID_EX_47), .IN2(ID_EX_46), .IN3(sp_en), .QN(n56) );
  AND4X1 U61 ( .IN1(n58), .IN2(n59), .IN3(wb_valid), .IN4(n60), .Q(n48) );
  XNOR2X1 U62 ( .IN1(ID_EX_46), .IN2(wb_rd[0]), .Q(n59) );
  XNOR2X1 U63 ( .IN1(ID_EX_47), .IN2(wb_rd[1]), .Q(n58) );
  XNOR2X1 U64 ( .IN1(ID_EX_47), .IN2(n6), .Q(n62) );
  XNOR2X1 U65 ( .IN1(ID_EX_46), .IN2(mem_rd[0]), .Q(n61) );
  AO221X1 U66 ( .IN1(ID_EX[7]), .IN2(n63), .IN3(n64), .IN4(sp_data[7]), .IN5(
        n65), .Q(s1_tmp[7]) );
  AO22X1 U67 ( .IN1(n66), .IN2(mem_data[7]), .IN3(n67), .IN4(wb_data[7]), .Q(
        n65) );
  AO221X1 U68 ( .IN1(ID_EX[6]), .IN2(n63), .IN3(n64), .IN4(sp_data[6]), .IN5(
        n68), .Q(s1_tmp[6]) );
  AO22X1 U69 ( .IN1(n66), .IN2(mem_data[6]), .IN3(n67), .IN4(wb_data[6]), .Q(
        n68) );
  AO221X1 U70 ( .IN1(ID_EX[5]), .IN2(n63), .IN3(n64), .IN4(sp_data[5]), .IN5(
        n69), .Q(s1_tmp[5]) );
  AO22X1 U71 ( .IN1(n66), .IN2(mem_data[5]), .IN3(n67), .IN4(wb_data[5]), .Q(
        n69) );
  AO221X1 U72 ( .IN1(ID_EX[4]), .IN2(n63), .IN3(n64), .IN4(sp_data[4]), .IN5(
        n70), .Q(s1_tmp[4]) );
  AO22X1 U73 ( .IN1(n66), .IN2(mem_data[4]), .IN3(n67), .IN4(wb_data[4]), .Q(
        n70) );
  AO221X1 U74 ( .IN1(ID_EX[3]), .IN2(n63), .IN3(n64), .IN4(sp_data[3]), .IN5(
        n71), .Q(s1_tmp[3]) );
  AO22X1 U75 ( .IN1(n66), .IN2(mem_data[3]), .IN3(n67), .IN4(wb_data[3]), .Q(
        n71) );
  AO221X1 U76 ( .IN1(ID_EX[2]), .IN2(n63), .IN3(n64), .IN4(sp_data[2]), .IN5(
        n72), .Q(s1_tmp[2]) );
  AO22X1 U77 ( .IN1(n66), .IN2(mem_data[2]), .IN3(n67), .IN4(wb_data[2]), .Q(
        n72) );
  AO221X1 U78 ( .IN1(ID_EX[1]), .IN2(n63), .IN3(n64), .IN4(sp_data[1]), .IN5(
        n73), .Q(s1_tmp[1]) );
  AO22X1 U79 ( .IN1(n66), .IN2(mem_data[1]), .IN3(n67), .IN4(wb_data[1]), .Q(
        n73) );
  AO221X1 U80 ( .IN1(ID_EX[0]), .IN2(n63), .IN3(n64), .IN4(sp_data[0]), .IN5(
        n74), .Q(s1_tmp[0]) );
  AO22X1 U81 ( .IN1(n66), .IN2(mem_data[0]), .IN3(n67), .IN4(wb_data[0]), .Q(
        n74) );
  AND2X1 U82 ( .IN1(n76), .IN2(n75), .Q(n63) );
  NAND4X0 U83 ( .IN1(ID_EX_40), .IN2(ID_EX[9]), .IN3(ID_EX[8]), .IN4(sp_en), 
        .QN(n75) );
  AND4X1 U84 ( .IN1(wb_valid), .IN2(n77), .IN3(ID_EX_40), .IN4(n78), .Q(n67)
         );
  XOR2X1 U85 ( .IN1(wb_rd[1]), .IN2(ID_EX[9]), .Q(n80) );
  XOR2X1 U86 ( .IN1(wb_rd[0]), .IN2(ID_EX[8]), .Q(n79) );
  AND3X1 U87 ( .IN1(ID_EX_40), .IN2(mem_valid), .IN3(n14), .Q(n66) );
  XNOR2X1 U89 ( .IN1(mem_rd[0]), .IN2(ID_EX[8]), .Q(n81) );
  AO22X1 U90 ( .IN1(CCR[3]), .IN2(n83), .IN3(flags_in[3]), .IN4(n17), .Q(
        flags_out[3]) );
  AO22X1 U91 ( .IN1(CCR[2]), .IN2(n16), .IN3(flags_in[2]), .IN4(n84), .Q(
        flags_out[2]) );
  OA21X1 U92 ( .IN1(n85), .IN2(n86), .IN3(n17), .Q(n84) );
  OA22X1 U93 ( .IN1(n20), .IN2(n87), .IN3(ID_EX[31]), .IN4(n18), .Q(n85) );
  AO22X1 U94 ( .IN1(CCR[1]), .IN2(n15), .IN3(flags_in[1]), .IN4(n88), .Q(
        flags_out[1]) );
  AO22X1 U95 ( .IN1(CCR[0]), .IN2(n15), .IN3(flags_in[0]), .IN4(n88), .Q(
        flags_out[0]) );
  OA21X1 U96 ( .IN1(n89), .IN2(n86), .IN3(n17), .Q(n88) );
  NOR3X0 U97 ( .IN1(n86), .IN2(ID_EX[30]), .IN3(n18), .QN(n83) );
  OA22X1 U98 ( .IN1(n19), .IN2(n90), .IN3(ID_EX[30]), .IN4(n20), .Q(n89) );
  AO222X1 U99 ( .IN1(n91), .IN2(ID_EX_43), .IN3(ID_EX_45), .IN4(n92), .IN5(n93), .IN6(n27), .Q(branch) );
  NAND3X0 U100 ( .IN1(flags_in[0]), .IN2(n25), .IN3(ID_EX_44), .QN(n95) );
  OAI21X1 U101 ( .IN1(n26), .IN2(flags_in[1]), .IN3(ID_EX_43), .QN(n94) );
  OA22X1 U102 ( .IN1(n26), .IN2(CCR[0]), .IN3(ID_EX_44), .IN4(n29), .Q(n96) );
  AND2X1 U103 ( .IN1(n26), .IN2(flags_in[3]), .Q(n91) );
  AO22X1 U104 ( .IN1(ID_EX_34), .IN2(ID_EX[27]), .IN3(EX_MEM[15]), .IN4(n21), 
        .Q(alu_b[7]) );
  AO22X1 U105 ( .IN1(ID_EX[26]), .IN2(ID_EX_34), .IN3(EX_MEM[14]), .IN4(n21), 
        .Q(alu_b[6]) );
  AO22X1 U106 ( .IN1(ID_EX[25]), .IN2(ID_EX_34), .IN3(EX_MEM[13]), .IN4(n21), 
        .Q(alu_b[5]) );
  AO22X1 U107 ( .IN1(ID_EX[24]), .IN2(ID_EX_34), .IN3(EX_MEM[12]), .IN4(n21), 
        .Q(alu_b[4]) );
  AO22X1 U108 ( .IN1(ID_EX[23]), .IN2(ID_EX_34), .IN3(EX_MEM[11]), .IN4(n21), 
        .Q(alu_b[3]) );
  AO22X1 U109 ( .IN1(ID_EX[22]), .IN2(ID_EX_34), .IN3(EX_MEM[10]), .IN4(n21), 
        .Q(alu_b[2]) );
  AO22X1 U110 ( .IN1(ID_EX[21]), .IN2(ID_EX_34), .IN3(EX_MEM[9]), .IN4(n21), 
        .Q(alu_b[1]) );
  AO22X1 U111 ( .IN1(ID_EX[20]), .IN2(ID_EX_34), .IN3(EX_MEM[8]), .IN4(n21), 
        .Q(alu_b[0]) );
  AO22X1 U113 ( .IN1(n100), .IN2(mem_data[1]), .IN3(n101), .IN4(wb_data[1]), 
        .Q(n99) );
  AO221X1 U114 ( .IN1(ID_EX[10]), .IN2(n97), .IN3(n98), .IN4(sp_data[0]), 
        .IN5(n102), .Q(EX_MEM[8]) );
  AO22X1 U115 ( .IN1(n100), .IN2(mem_data[0]), .IN3(n101), .IN4(wb_data[0]), 
        .Q(n102) );
  AO22X1 U116 ( .IN1(result[7]), .IN2(n103), .IN3(IN_PORT[7]), .IN4(n22), .Q(
        EX_MEM[7]) );
  AO22X1 U117 ( .IN1(result[6]), .IN2(n103), .IN3(IN_PORT[6]), .IN4(n22), .Q(
        EX_MEM[6]) );
  AO22X1 U118 ( .IN1(result[5]), .IN2(n103), .IN3(IN_PORT[5]), .IN4(n22), .Q(
        EX_MEM[5]) );
  AO22X1 U119 ( .IN1(result[4]), .IN2(n103), .IN3(IN_PORT[4]), .IN4(n22), .Q(
        EX_MEM[4]) );
  AO22X1 U120 ( .IN1(result[3]), .IN2(n103), .IN3(IN_PORT[3]), .IN4(n22), .Q(
        EX_MEM[3]) );
  AO22X1 U121 ( .IN1(result[2]), .IN2(n103), .IN3(IN_PORT[2]), .IN4(n22), .Q(
        EX_MEM[2]) );
  AND4X1 U122 ( .IN1(mem_acc_mode[0]), .IN2(ID_EX_38), .IN3(n104), .IN4(n31), 
        .Q(N120) );
  NAND3X0 U123 ( .IN1(n107), .IN2(ID_EX_41), .IN3(n108), .QN(n106) );
  XNOR2X1 U124 ( .IN1(stall_Rd[0]), .IN2(ID_EX[18]), .Q(n108) );
  XNOR2X1 U125 ( .IN1(stall_Rd[1]), .IN2(ID_EX[19]), .Q(n107) );
  NAND3X0 U126 ( .IN1(n109), .IN2(ID_EX_40), .IN3(n110), .QN(n105) );
  XNOR2X1 U127 ( .IN1(stall_Rd[0]), .IN2(ID_EX[8]), .Q(n110) );
  XNOR2X1 U128 ( .IN1(stall_Rd[1]), .IN2(ID_EX[9]), .Q(n109) );
  AO22X1 U129 ( .IN1(result[1]), .IN2(n103), .IN3(IN_PORT[1]), .IN4(n22), .Q(
        EX_MEM[1]) );
  AO221X1 U130 ( .IN1(ID_EX[17]), .IN2(n3), .IN3(n10), .IN4(sp_data[7]), .IN5(
        n111), .Q(EX_MEM[15]) );
  AO221X1 U132 ( .IN1(ID_EX[16]), .IN2(n3), .IN3(n10), .IN4(sp_data[6]), .IN5(
        n112), .Q(EX_MEM[14]) );
  AO22X1 U133 ( .IN1(n100), .IN2(mem_data[6]), .IN3(n101), .IN4(wb_data[6]), 
        .Q(n112) );
  AO221X1 U134 ( .IN1(ID_EX[15]), .IN2(n3), .IN3(n10), .IN4(sp_data[5]), .IN5(
        n113), .Q(EX_MEM[13]) );
  AO22X1 U135 ( .IN1(n100), .IN2(mem_data[5]), .IN3(n101), .IN4(wb_data[5]), 
        .Q(n113) );
  AO221X1 U136 ( .IN1(ID_EX[14]), .IN2(n3), .IN3(n10), .IN4(sp_data[4]), .IN5(
        n114), .Q(EX_MEM[12]) );
  AO22X1 U137 ( .IN1(n100), .IN2(mem_data[4]), .IN3(n101), .IN4(wb_data[4]), 
        .Q(n114) );
  AO221X1 U138 ( .IN1(ID_EX[13]), .IN2(n3), .IN3(n10), .IN4(sp_data[3]), .IN5(
        n115), .Q(EX_MEM[11]) );
  AO22X1 U139 ( .IN1(n100), .IN2(mem_data[3]), .IN3(n101), .IN4(wb_data[3]), 
        .Q(n115) );
  AO22X1 U141 ( .IN1(n100), .IN2(mem_data[2]), .IN3(n101), .IN4(wb_data[2]), 
        .Q(n116) );
  NAND4X0 U143 ( .IN1(ID_EX_41), .IN2(ID_EX[19]), .IN3(ID_EX[18]), .IN4(sp_en), 
        .QN(n117) );
  XOR2X1 U145 ( .IN1(wb_rd[1]), .IN2(ID_EX[19]), .Q(n122) );
  XOR2X1 U146 ( .IN1(wb_rd[0]), .IN2(ID_EX[18]), .Q(n121) );
  XNOR2X1 U148 ( .IN1(mem_rd[1]), .IN2(ID_EX[19]), .Q(n124) );
  XNOR2X1 U149 ( .IN1(mem_rd[0]), .IN2(ID_EX[18]), .Q(n123) );
  AO22X1 U150 ( .IN1(result[0]), .IN2(n103), .IN3(IN_PORT[0]), .IN4(n22), .Q(
        EX_MEM[0]) );
  NAND3X0 U151 ( .IN1(\ID_EX[36] ), .IN2(n23), .IN3(\ID_EX[37] ), .QN(n103) );
  ALSU alu0 ( .a(s1_tmp), .b(alu_b), .s(ID_EX[31:28]), .cin(flags_in[2]), .F(
        result), .cout(CCR[2]), .zero(CCR[0]), .negative(CCR[1]), .overflow(
        CCR[3]) );
  XNOR2X1 U3 ( .IN1(mem_rd[1]), .IN2(ID_EX[9]), .Q(n82) );
  NBUFFX2 U4 ( .IN(mem_rd[1]), .Q(n6) );
  INVX0 U5 ( .IN(n117), .QN(n5) );
  INVX0 U6 ( .IN(n2), .QN(n9) );
  NBUFFX2 U7 ( .IN(n97), .Q(n1) );
  AO221X1 U8 ( .IN1(ID_EX[12]), .IN2(n1), .IN3(n2), .IN4(sp_data[2]), .IN5(
        n116), .Q(EX_MEM[10]) );
  AO221X1 U9 ( .IN1(ID_EX[11]), .IN2(n97), .IN3(n2), .IN4(sp_data[1]), .IN5(
        n99), .Q(EX_MEM[9]) );
  NOR2X0 U10 ( .IN1(n7), .IN2(n117), .QN(n2) );
  NOR2X0 U11 ( .IN1(n7), .IN2(n117), .QN(n98) );
  NBUFFX2 U12 ( .IN(n1), .Q(n3) );
  NOR2X0 U13 ( .IN1(n100), .IN2(n4), .QN(n97) );
  OR2X1 U14 ( .IN1(n101), .IN2(n5), .Q(n4) );
  OR2X1 U15 ( .IN1(n100), .IN2(n101), .Q(n7) );
  AND3X2 U16 ( .IN1(n8), .IN2(mem_valid), .IN3(ID_EX_41), .Q(n100) );
  AND2X1 U17 ( .IN1(n123), .IN2(n124), .Q(n8) );
  NOR2X1 U18 ( .IN1(n75), .IN2(n13), .QN(n64) );
  INVX0 U19 ( .IN(n9), .QN(n10) );
  INVX0 U20 ( .IN(n76), .QN(n13) );
  NOR2X0 U21 ( .IN1(n66), .IN2(n67), .QN(n76) );
  NOR2X0 U22 ( .IN1(n30), .IN2(n60), .QN(n47) );
  INVX0 U23 ( .IN(mem_valid), .QN(n30) );
  NOR2X0 U24 ( .IN1(n56), .IN2(n28), .QN(n45) );
  INVX0 U25 ( .IN(n57), .QN(n28) );
  NOR2X0 U26 ( .IN1(n47), .IN2(n48), .QN(n57) );
  INVX0 U27 ( .IN(n83), .QN(n17) );
  INVX0 U28 ( .IN(n88), .QN(n15) );
  INVX0 U29 ( .IN(n103), .QN(n22) );
  NOR2X0 U30 ( .IN1(n79), .IN2(n80), .QN(n78) );
  INVX0 U31 ( .IN(n77), .QN(n14) );
  INVX0 U32 ( .IN(ID_EX_45), .QN(n27) );
  NAND2X0 U33 ( .IN1(n94), .IN2(n95), .QN(n93) );
  NOR2X0 U34 ( .IN1(n121), .IN2(n122), .QN(n120) );
  INVX0 U35 ( .IN(flags_in[2]), .QN(n29) );
  INVX0 U36 ( .IN(n84), .QN(n16) );
  NAND2X0 U37 ( .IN1(n123), .IN2(n124), .QN(n119) );
  NAND2X0 U38 ( .IN1(n81), .IN2(n82), .QN(n77) );
  INVX0 U39 ( .IN(ID_EX_34), .QN(n21) );
  INVX0 U40 ( .IN(mem_acc_mode[2]), .QN(n31) );
  NAND2X0 U41 ( .IN1(n105), .IN2(n106), .QN(n104) );
  NAND2X0 U42 ( .IN1(n61), .IN2(n62), .QN(n60) );
  INVX0 U88 ( .IN(ID_EX_43), .QN(n25) );
  INVX0 U112 ( .IN(ID_EX[29]), .QN(n18) );
  INVX0 U131 ( .IN(ID_EX[31]), .QN(n20) );
  INVX0 U140 ( .IN(ID_EX[30]), .QN(n19) );
  NAND2X0 U142 ( .IN1(n18), .IN2(n20), .QN(n90) );
  NAND2X0 U144 ( .IN1(ID_EX[30]), .IN2(n18), .QN(n87) );
  NAND2X0 U147 ( .IN1(ID_EX_39), .IN2(ID_EX_38), .QN(n86) );
  INVX0 U152 ( .IN(ID_EX_44), .QN(n26) );
  INVX0 U153 ( .IN(\ID_EX[35] ), .QN(n23) );
  NOR2X0 U154 ( .IN1(N120), .IN2(n24), .QN(EX_MEM[21]) );
  INVX0 U155 ( .IN(ID_EX_38), .QN(n24) );
  NAND2X0 U156 ( .IN1(n100), .IN2(mem_data[7]), .QN(n11) );
  NAND2X0 U157 ( .IN1(n101), .IN2(wb_data[7]), .QN(n12) );
  NAND2X0 U158 ( .IN1(n12), .IN2(n11), .QN(n111) );
  AND4X2 U159 ( .IN1(n119), .IN2(wb_valid), .IN3(ID_EX_41), .IN4(n120), .Q(
        n101) );
  NOR2X0 U160 ( .IN1(n96), .IN2(ID_EX_43), .QN(n92) );
endmodule


module my_DFF_1_100 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_99 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_98 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_97 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_nDFF_n4 ( clk, rst, e, d, q );
  input [3:0] d;
  output [3:0] q;
  input clk, rst, e;


  my_DFF_1_100 fx_0 ( .d(d[0]), .clk(clk), .rst(rst), .e(e), .q(q[0]) );
  my_DFF_1_99 fx_1 ( .d(d[1]), .clk(clk), .rst(rst), .e(e), .q(q[1]) );
  my_DFF_1_98 fx_2 ( .d(d[2]), .clk(clk), .rst(rst), .e(e), .q(q[2]) );
  my_DFF_1_97 fx_3 ( .d(d[3]), .clk(clk), .rst(rst), .e(e), .q(q[3]) );
endmodule


module my_DFF_1_96 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_95 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_94 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_93 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_92 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_91 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_90 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_89 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_88 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_87 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_86 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_85 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_84 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_83 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_82 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_81 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_80 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_79 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_78 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n7, n1, n4, n5, n6;

  DFFARX1 q_reg ( .D(n6), .CLK(clk), .RSTB(n4), .Q(n7), .QN(n1) );
  AO22X1 U3 ( .IN1(n7), .IN2(n5), .IN3(e), .IN4(d), .Q(n6) );
  INVX0 U2 ( .IN(rst), .QN(n4) );
  INVX0 U4 ( .IN(e), .QN(n5) );
  INVX0 U5 ( .IN(n1), .QN(q) );
endmodule


module my_DFF_1_77 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n7, n1, n4, n5, n6;

  DFFARX1 q_reg ( .D(n6), .CLK(clk), .RSTB(n4), .Q(n7), .QN(n1) );
  AO22X1 U3 ( .IN1(n7), .IN2(n5), .IN3(e), .IN4(d), .Q(n6) );
  INVX0 U2 ( .IN(rst), .QN(n4) );
  INVX0 U4 ( .IN(e), .QN(n5) );
  INVX0 U5 ( .IN(n1), .QN(q) );
endmodule


module my_DFF_1_76 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n7, n1, n4, n5, n6;

  DFFARX1 q_reg ( .D(n6), .CLK(clk), .RSTB(n4), .Q(n7), .QN(n1) );
  AO22X1 U3 ( .IN1(n7), .IN2(n5), .IN3(e), .IN4(d), .Q(n6) );
  INVX0 U2 ( .IN(n1), .QN(q) );
  INVX0 U4 ( .IN(rst), .QN(n4) );
  INVX0 U5 ( .IN(e), .QN(n5) );
endmodule


module my_DFF_1_75 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n7, n1, n4, n5, n6;

  DFFARX1 q_reg ( .D(n6), .CLK(clk), .RSTB(n4), .Q(n7), .QN(n1) );
  AO22X1 U3 ( .IN1(n7), .IN2(n5), .IN3(e), .IN4(d), .Q(n6) );
  INVX1 U2 ( .IN(n1), .QN(q) );
  INVX0 U4 ( .IN(rst), .QN(n4) );
  INVX0 U5 ( .IN(e), .QN(n5) );
endmodule


module my_DFF_1_74 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_73 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_72 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_71 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_70 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_69 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_68 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_67 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_66 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_65 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_nDFF_n32_2 ( clk, rst, e, d, q );
  input [31:0] d;
  output [31:0] q;
  input clk, rst, e;
  wire   n1, n2, n3;

  my_DFF_1_96 fx_0 ( .d(d[0]), .clk(clk), .rst(n3), .e(e), .q(q[0]) );
  my_DFF_1_95 fx_1 ( .d(d[1]), .clk(clk), .rst(n3), .e(e), .q(q[1]) );
  my_DFF_1_94 fx_2 ( .d(d[2]), .clk(clk), .rst(n3), .e(e), .q(q[2]) );
  my_DFF_1_93 fx_3 ( .d(d[3]), .clk(clk), .rst(n3), .e(e), .q(q[3]) );
  my_DFF_1_92 fx_4 ( .d(d[4]), .clk(clk), .rst(n3), .e(e), .q(q[4]) );
  my_DFF_1_91 fx_5 ( .d(d[5]), .clk(clk), .rst(n3), .e(e), .q(q[5]) );
  my_DFF_1_90 fx_6 ( .d(d[6]), .clk(clk), .rst(n3), .e(e), .q(q[6]) );
  my_DFF_1_89 fx_7 ( .d(d[7]), .clk(clk), .rst(n3), .e(e), .q(q[7]) );
  my_DFF_1_88 fx_8 ( .d(d[8]), .clk(clk), .rst(n2), .e(e), .q(q[8]) );
  my_DFF_1_87 fx_9 ( .d(d[9]), .clk(clk), .rst(n2), .e(e), .q(q[9]) );
  my_DFF_1_86 fx_10 ( .d(d[10]), .clk(clk), .rst(n2), .e(e), .q(q[10]) );
  my_DFF_1_85 fx_11 ( .d(d[11]), .clk(clk), .rst(n2), .e(e), .q(q[11]) );
  my_DFF_1_84 fx_12 ( .d(d[12]), .clk(clk), .rst(n2), .e(e), .q(q[12]) );
  my_DFF_1_83 fx_13 ( .d(d[13]), .clk(clk), .rst(n2), .e(e), .q(q[13]) );
  my_DFF_1_82 fx_14 ( .d(d[14]), .clk(clk), .rst(n2), .e(e), .q(q[14]) );
  my_DFF_1_81 fx_15 ( .d(d[15]), .clk(clk), .rst(n2), .e(e), .q(q[15]) );
  my_DFF_1_80 fx_16 ( .d(d[16]), .clk(clk), .rst(n2), .e(e), .q(q[16]) );
  my_DFF_1_79 fx_17 ( .d(d[17]), .clk(clk), .rst(n2), .e(e), .q(q[17]) );
  my_DFF_1_78 fx_18 ( .d(d[18]), .clk(clk), .rst(n2), .e(e), .q(q[18]) );
  my_DFF_1_77 fx_19 ( .d(d[19]), .clk(clk), .rst(n2), .e(e), .q(q[19]) );
  my_DFF_1_76 fx_20 ( .d(d[20]), .clk(clk), .rst(n1), .e(e), .q(q[20]) );
  my_DFF_1_75 fx_21 ( .d(d[21]), .clk(clk), .rst(n1), .e(e), .q(q[21]) );
  my_DFF_1_74 fx_22 ( .d(d[22]), .clk(clk), .rst(n1), .e(e), .q(q[22]) );
  my_DFF_1_73 fx_23 ( .d(d[23]), .clk(clk), .rst(n1), .e(e), .q(q[23]) );
  my_DFF_1_72 fx_24 ( .d(d[24]), .clk(clk), .rst(n1), .e(e), .q(q[24]) );
  my_DFF_1_71 fx_25 ( .d(d[25]), .clk(clk), .rst(n1), .e(e), .q(q[25]) );
  my_DFF_1_70 fx_26 ( .d(d[26]), .clk(clk), .rst(n1), .e(e), .q(q[26]) );
  my_DFF_1_69 fx_27 ( .d(d[27]), .clk(clk), .rst(n1), .e(e), .q(q[27]) );
  my_DFF_1_68 fx_28 ( .d(d[28]), .clk(clk), .rst(n1), .e(e), .q(q[28]) );
  my_DFF_1_67 fx_29 ( .d(d[29]), .clk(clk), .rst(n1), .e(e), .q(q[29]) );
  my_DFF_1_66 fx_30 ( .d(d[30]), .clk(clk), .rst(n1), .e(e), .q(q[30]) );
  my_DFF_1_65 fx_31 ( .d(d[31]), .clk(clk), .rst(n1), .e(e), .q(q[31]) );
  NBUFFX2 U1 ( .IN(rst), .Q(n2) );
  NBUFFX2 U2 ( .IN(rst), .Q(n1) );
  NBUFFX2 U3 ( .IN(rst), .Q(n3) );
endmodule


module data_ram_1 ( clk, R, W, address, datain, dataout, MFC );
  input [7:0] address;
  input [7:0] datain;
  output [7:0] dataout;
  input clk, R, W;
  output MFC;
  wire   \ram[0][7] , \ram[0][6] , \ram[0][5] , \ram[0][4] , \ram[0][3] ,
         \ram[0][2] , \ram[0][1] , \ram[0][0] , \ram[1][7] , \ram[1][6] ,
         \ram[1][5] , \ram[1][4] , \ram[1][3] , \ram[1][2] , \ram[1][1] ,
         \ram[1][0] , \ram[2][7] , \ram[2][6] , \ram[2][5] , \ram[2][4] ,
         \ram[2][3] , \ram[2][2] , \ram[2][1] , \ram[2][0] , \ram[3][7] ,
         \ram[3][6] , \ram[3][5] , \ram[3][4] , \ram[3][3] , \ram[3][2] ,
         \ram[3][1] , \ram[3][0] , \ram[4][7] , \ram[4][6] , \ram[4][5] ,
         \ram[4][4] , \ram[4][3] , \ram[4][2] , \ram[4][1] , \ram[4][0] ,
         \ram[5][7] , \ram[5][6] , \ram[5][5] , \ram[5][4] , \ram[5][3] ,
         \ram[5][2] , \ram[5][1] , \ram[5][0] , \ram[6][7] , \ram[6][6] ,
         \ram[6][5] , \ram[6][4] , \ram[6][3] , \ram[6][2] , \ram[6][1] ,
         \ram[6][0] , \ram[7][7] , \ram[7][6] , \ram[7][5] , \ram[7][4] ,
         \ram[7][3] , \ram[7][2] , \ram[7][1] , \ram[7][0] , \ram[8][7] ,
         \ram[8][6] , \ram[8][5] , \ram[8][4] , \ram[8][3] , \ram[8][2] ,
         \ram[8][1] , \ram[8][0] , \ram[9][7] , \ram[9][6] , \ram[9][5] ,
         \ram[9][4] , \ram[9][3] , \ram[9][2] , \ram[9][1] , \ram[9][0] ,
         \ram[10][7] , \ram[10][6] , \ram[10][5] , \ram[10][4] , \ram[10][3] ,
         \ram[10][2] , \ram[10][1] , \ram[10][0] , \ram[11][7] , \ram[11][6] ,
         \ram[11][5] , \ram[11][4] , \ram[11][3] , \ram[11][2] , \ram[11][1] ,
         \ram[11][0] , \ram[12][7] , \ram[12][6] , \ram[12][5] , \ram[12][4] ,
         \ram[12][3] , \ram[12][2] , \ram[12][1] , \ram[12][0] , \ram[13][7] ,
         \ram[13][6] , \ram[13][5] , \ram[13][4] , \ram[13][3] , \ram[13][2] ,
         \ram[13][1] , \ram[13][0] , \ram[14][7] , \ram[14][6] , \ram[14][5] ,
         \ram[14][4] , \ram[14][3] , \ram[14][2] , \ram[14][1] , \ram[14][0] ,
         \ram[15][7] , \ram[15][6] , \ram[15][5] , \ram[15][4] , \ram[15][3] ,
         \ram[15][2] , \ram[15][1] , \ram[15][0] , \ram[16][7] , \ram[16][6] ,
         \ram[16][5] , \ram[16][4] , \ram[16][3] , \ram[16][2] , \ram[16][1] ,
         \ram[16][0] , \ram[17][7] , \ram[17][6] , \ram[17][5] , \ram[17][4] ,
         \ram[17][3] , \ram[17][2] , \ram[17][1] , \ram[17][0] , \ram[18][7] ,
         \ram[18][6] , \ram[18][5] , \ram[18][4] , \ram[18][3] , \ram[18][2] ,
         \ram[18][1] , \ram[18][0] , \ram[19][7] , \ram[19][6] , \ram[19][5] ,
         \ram[19][4] , \ram[19][3] , \ram[19][2] , \ram[19][1] , \ram[19][0] ,
         \ram[20][7] , \ram[20][6] , \ram[20][5] , \ram[20][4] , \ram[20][3] ,
         \ram[20][2] , \ram[20][1] , \ram[20][0] , \ram[21][7] , \ram[21][6] ,
         \ram[21][5] , \ram[21][4] , \ram[21][3] , \ram[21][2] , \ram[21][1] ,
         \ram[21][0] , \ram[22][7] , \ram[22][6] , \ram[22][5] , \ram[22][4] ,
         \ram[22][3] , \ram[22][2] , \ram[22][1] , \ram[22][0] , \ram[23][7] ,
         \ram[23][6] , \ram[23][5] , \ram[23][4] , \ram[23][3] , \ram[23][2] ,
         \ram[23][1] , \ram[23][0] , \ram[24][7] , \ram[24][6] , \ram[24][5] ,
         \ram[24][4] , \ram[24][3] , \ram[24][2] , \ram[24][1] , \ram[24][0] ,
         \ram[25][7] , \ram[25][6] , \ram[25][5] , \ram[25][4] , \ram[25][3] ,
         \ram[25][2] , \ram[25][1] , \ram[25][0] , \ram[26][7] , \ram[26][6] ,
         \ram[26][5] , \ram[26][4] , \ram[26][3] , \ram[26][2] , \ram[26][1] ,
         \ram[26][0] , \ram[27][7] , \ram[27][6] , \ram[27][5] , \ram[27][4] ,
         \ram[27][3] , \ram[27][2] , \ram[27][1] , \ram[27][0] , \ram[28][7] ,
         \ram[28][6] , \ram[28][5] , \ram[28][4] , \ram[28][3] , \ram[28][2] ,
         \ram[28][1] , \ram[28][0] , \ram[29][7] , \ram[29][6] , \ram[29][5] ,
         \ram[29][4] , \ram[29][3] , \ram[29][2] , \ram[29][1] , \ram[29][0] ,
         \ram[30][7] , \ram[30][6] , \ram[30][5] , \ram[30][4] , \ram[30][3] ,
         \ram[30][2] , \ram[30][1] , \ram[30][0] , \ram[31][7] , \ram[31][6] ,
         \ram[31][5] , \ram[31][4] , \ram[31][3] , \ram[31][2] , \ram[31][1] ,
         \ram[31][0] , \ram[32][7] , \ram[32][6] , \ram[32][5] , \ram[32][4] ,
         \ram[32][3] , \ram[32][2] , \ram[32][1] , \ram[32][0] , \ram[33][7] ,
         \ram[33][6] , \ram[33][5] , \ram[33][4] , \ram[33][3] , \ram[33][2] ,
         \ram[33][1] , \ram[33][0] , \ram[34][7] , \ram[34][6] , \ram[34][5] ,
         \ram[34][4] , \ram[34][3] , \ram[34][2] , \ram[34][1] , \ram[34][0] ,
         \ram[35][7] , \ram[35][6] , \ram[35][5] , \ram[35][4] , \ram[35][3] ,
         \ram[35][2] , \ram[35][1] , \ram[35][0] , \ram[36][7] , \ram[36][6] ,
         \ram[36][5] , \ram[36][4] , \ram[36][3] , \ram[36][2] , \ram[36][1] ,
         \ram[36][0] , \ram[37][7] , \ram[37][6] , \ram[37][5] , \ram[37][4] ,
         \ram[37][3] , \ram[37][2] , \ram[37][1] , \ram[37][0] , \ram[38][7] ,
         \ram[38][6] , \ram[38][5] , \ram[38][4] , \ram[38][3] , \ram[38][2] ,
         \ram[38][1] , \ram[38][0] , \ram[39][7] , \ram[39][6] , \ram[39][5] ,
         \ram[39][4] , \ram[39][3] , \ram[39][2] , \ram[39][1] , \ram[39][0] ,
         \ram[40][7] , \ram[40][6] , \ram[40][5] , \ram[40][4] , \ram[40][3] ,
         \ram[40][2] , \ram[40][1] , \ram[40][0] , \ram[41][7] , \ram[41][6] ,
         \ram[41][5] , \ram[41][4] , \ram[41][3] , \ram[41][2] , \ram[41][1] ,
         \ram[41][0] , \ram[42][7] , \ram[42][6] , \ram[42][5] , \ram[42][4] ,
         \ram[42][3] , \ram[42][2] , \ram[42][1] , \ram[42][0] , \ram[43][7] ,
         \ram[43][6] , \ram[43][5] , \ram[43][4] , \ram[43][3] , \ram[43][2] ,
         \ram[43][1] , \ram[43][0] , \ram[44][7] , \ram[44][6] , \ram[44][5] ,
         \ram[44][4] , \ram[44][3] , \ram[44][2] , \ram[44][1] , \ram[44][0] ,
         \ram[45][7] , \ram[45][6] , \ram[45][5] , \ram[45][4] , \ram[45][3] ,
         \ram[45][2] , \ram[45][1] , \ram[45][0] , \ram[46][7] , \ram[46][6] ,
         \ram[46][5] , \ram[46][4] , \ram[46][3] , \ram[46][2] , \ram[46][1] ,
         \ram[46][0] , \ram[47][7] , \ram[47][6] , \ram[47][5] , \ram[47][4] ,
         \ram[47][3] , \ram[47][2] , \ram[47][1] , \ram[47][0] , \ram[48][7] ,
         \ram[48][6] , \ram[48][5] , \ram[48][4] , \ram[48][3] , \ram[48][2] ,
         \ram[48][1] , \ram[48][0] , \ram[49][7] , \ram[49][6] , \ram[49][5] ,
         \ram[49][4] , \ram[49][3] , \ram[49][2] , \ram[49][1] , \ram[49][0] ,
         \ram[50][7] , \ram[50][6] , \ram[50][5] , \ram[50][4] , \ram[50][3] ,
         \ram[50][2] , \ram[50][1] , \ram[50][0] , \ram[51][7] , \ram[51][6] ,
         \ram[51][5] , \ram[51][4] , \ram[51][3] , \ram[51][2] , \ram[51][1] ,
         \ram[51][0] , \ram[52][7] , \ram[52][6] , \ram[52][5] , \ram[52][4] ,
         \ram[52][3] , \ram[52][2] , \ram[52][1] , \ram[52][0] , \ram[53][7] ,
         \ram[53][6] , \ram[53][5] , \ram[53][4] , \ram[53][3] , \ram[53][2] ,
         \ram[53][1] , \ram[53][0] , \ram[54][7] , \ram[54][6] , \ram[54][5] ,
         \ram[54][4] , \ram[54][3] , \ram[54][2] , \ram[54][1] , \ram[54][0] ,
         \ram[55][7] , \ram[55][6] , \ram[55][5] , \ram[55][4] , \ram[55][3] ,
         \ram[55][2] , \ram[55][1] , \ram[55][0] , \ram[56][7] , \ram[56][6] ,
         \ram[56][5] , \ram[56][4] , \ram[56][3] , \ram[56][2] , \ram[56][1] ,
         \ram[56][0] , \ram[57][7] , \ram[57][6] , \ram[57][5] , \ram[57][4] ,
         \ram[57][3] , \ram[57][2] , \ram[57][1] , \ram[57][0] , \ram[58][7] ,
         \ram[58][6] , \ram[58][5] , \ram[58][4] , \ram[58][3] , \ram[58][2] ,
         \ram[58][1] , \ram[58][0] , \ram[59][7] , \ram[59][6] , \ram[59][5] ,
         \ram[59][4] , \ram[59][3] , \ram[59][2] , \ram[59][1] , \ram[59][0] ,
         \ram[60][7] , \ram[60][6] , \ram[60][5] , \ram[60][4] , \ram[60][3] ,
         \ram[60][2] , \ram[60][1] , \ram[60][0] , \ram[61][7] , \ram[61][6] ,
         \ram[61][5] , \ram[61][4] , \ram[61][3] , \ram[61][2] , \ram[61][1] ,
         \ram[61][0] , \ram[62][7] , \ram[62][6] , \ram[62][5] , \ram[62][4] ,
         \ram[62][3] , \ram[62][2] , \ram[62][1] , \ram[62][0] , \ram[63][7] ,
         \ram[63][6] , \ram[63][5] , \ram[63][4] , \ram[63][3] , \ram[63][2] ,
         \ram[63][1] , \ram[63][0] , \ram[64][7] , \ram[64][6] , \ram[64][5] ,
         \ram[64][4] , \ram[64][3] , \ram[64][2] , \ram[64][1] , \ram[64][0] ,
         \ram[65][7] , \ram[65][6] , \ram[65][5] , \ram[65][4] , \ram[65][3] ,
         \ram[65][2] , \ram[65][1] , \ram[65][0] , \ram[66][7] , \ram[66][6] ,
         \ram[66][5] , \ram[66][4] , \ram[66][3] , \ram[66][2] , \ram[66][1] ,
         \ram[66][0] , \ram[67][7] , \ram[67][6] , \ram[67][5] , \ram[67][4] ,
         \ram[67][3] , \ram[67][2] , \ram[67][1] , \ram[67][0] , \ram[68][7] ,
         \ram[68][6] , \ram[68][5] , \ram[68][4] , \ram[68][3] , \ram[68][2] ,
         \ram[68][1] , \ram[68][0] , \ram[69][7] , \ram[69][6] , \ram[69][5] ,
         \ram[69][4] , \ram[69][3] , \ram[69][2] , \ram[69][1] , \ram[69][0] ,
         \ram[70][7] , \ram[70][6] , \ram[70][5] , \ram[70][4] , \ram[70][3] ,
         \ram[70][2] , \ram[70][1] , \ram[70][0] , \ram[71][7] , \ram[71][6] ,
         \ram[71][5] , \ram[71][4] , \ram[71][3] , \ram[71][2] , \ram[71][1] ,
         \ram[71][0] , \ram[72][7] , \ram[72][6] , \ram[72][5] , \ram[72][4] ,
         \ram[72][3] , \ram[72][2] , \ram[72][1] , \ram[72][0] , \ram[73][7] ,
         \ram[73][6] , \ram[73][5] , \ram[73][4] , \ram[73][3] , \ram[73][2] ,
         \ram[73][1] , \ram[73][0] , \ram[74][7] , \ram[74][6] , \ram[74][5] ,
         \ram[74][4] , \ram[74][3] , \ram[74][2] , \ram[74][1] , \ram[74][0] ,
         \ram[75][7] , \ram[75][6] , \ram[75][5] , \ram[75][4] , \ram[75][3] ,
         \ram[75][2] , \ram[75][1] , \ram[75][0] , \ram[76][7] , \ram[76][6] ,
         \ram[76][5] , \ram[76][4] , \ram[76][3] , \ram[76][2] , \ram[76][1] ,
         \ram[76][0] , \ram[77][7] , \ram[77][6] , \ram[77][5] , \ram[77][4] ,
         \ram[77][3] , \ram[77][2] , \ram[77][1] , \ram[77][0] , \ram[78][7] ,
         \ram[78][6] , \ram[78][5] , \ram[78][4] , \ram[78][3] , \ram[78][2] ,
         \ram[78][1] , \ram[78][0] , \ram[79][7] , \ram[79][6] , \ram[79][5] ,
         \ram[79][4] , \ram[79][3] , \ram[79][2] , \ram[79][1] , \ram[79][0] ,
         \ram[80][7] , \ram[80][6] , \ram[80][5] , \ram[80][4] , \ram[80][3] ,
         \ram[80][2] , \ram[80][1] , \ram[80][0] , \ram[81][7] , \ram[81][6] ,
         \ram[81][5] , \ram[81][4] , \ram[81][3] , \ram[81][2] , \ram[81][1] ,
         \ram[81][0] , \ram[82][7] , \ram[82][6] , \ram[82][5] , \ram[82][4] ,
         \ram[82][3] , \ram[82][2] , \ram[82][1] , \ram[82][0] , \ram[83][7] ,
         \ram[83][6] , \ram[83][5] , \ram[83][4] , \ram[83][3] , \ram[83][2] ,
         \ram[83][1] , \ram[83][0] , \ram[84][7] , \ram[84][6] , \ram[84][5] ,
         \ram[84][4] , \ram[84][3] , \ram[84][2] , \ram[84][1] , \ram[84][0] ,
         \ram[85][7] , \ram[85][6] , \ram[85][5] , \ram[85][4] , \ram[85][3] ,
         \ram[85][2] , \ram[85][1] , \ram[85][0] , \ram[86][7] , \ram[86][6] ,
         \ram[86][5] , \ram[86][4] , \ram[86][3] , \ram[86][2] , \ram[86][1] ,
         \ram[86][0] , \ram[87][7] , \ram[87][6] , \ram[87][5] , \ram[87][4] ,
         \ram[87][3] , \ram[87][2] , \ram[87][1] , \ram[87][0] , \ram[88][7] ,
         \ram[88][6] , \ram[88][5] , \ram[88][4] , \ram[88][3] , \ram[88][2] ,
         \ram[88][1] , \ram[88][0] , \ram[89][7] , \ram[89][6] , \ram[89][5] ,
         \ram[89][4] , \ram[89][3] , \ram[89][2] , \ram[89][1] , \ram[89][0] ,
         \ram[90][7] , \ram[90][6] , \ram[90][5] , \ram[90][4] , \ram[90][3] ,
         \ram[90][2] , \ram[90][1] , \ram[90][0] , \ram[91][7] , \ram[91][6] ,
         \ram[91][5] , \ram[91][4] , \ram[91][3] , \ram[91][2] , \ram[91][1] ,
         \ram[91][0] , \ram[92][7] , \ram[92][6] , \ram[92][5] , \ram[92][4] ,
         \ram[92][3] , \ram[92][2] , \ram[92][1] , \ram[92][0] , \ram[93][7] ,
         \ram[93][6] , \ram[93][5] , \ram[93][4] , \ram[93][3] , \ram[93][2] ,
         \ram[93][1] , \ram[93][0] , \ram[94][7] , \ram[94][6] , \ram[94][5] ,
         \ram[94][4] , \ram[94][3] , \ram[94][2] , \ram[94][1] , \ram[94][0] ,
         \ram[95][7] , \ram[95][6] , \ram[95][5] , \ram[95][4] , \ram[95][3] ,
         \ram[95][2] , \ram[95][1] , \ram[95][0] , \ram[96][7] , \ram[96][6] ,
         \ram[96][5] , \ram[96][4] , \ram[96][3] , \ram[96][2] , \ram[96][1] ,
         \ram[96][0] , \ram[97][7] , \ram[97][6] , \ram[97][5] , \ram[97][4] ,
         \ram[97][3] , \ram[97][2] , \ram[97][1] , \ram[97][0] , \ram[98][7] ,
         \ram[98][6] , \ram[98][5] , \ram[98][4] , \ram[98][3] , \ram[98][2] ,
         \ram[98][1] , \ram[98][0] , \ram[99][7] , \ram[99][6] , \ram[99][5] ,
         \ram[99][4] , \ram[99][3] , \ram[99][2] , \ram[99][1] , \ram[99][0] ,
         \ram[100][7] , \ram[100][6] , \ram[100][5] , \ram[100][4] ,
         \ram[100][3] , \ram[100][2] , \ram[100][1] , \ram[100][0] ,
         \ram[101][7] , \ram[101][6] , \ram[101][5] , \ram[101][4] ,
         \ram[101][3] , \ram[101][2] , \ram[101][1] , \ram[101][0] ,
         \ram[102][7] , \ram[102][6] , \ram[102][5] , \ram[102][4] ,
         \ram[102][3] , \ram[102][2] , \ram[102][1] , \ram[102][0] ,
         \ram[103][7] , \ram[103][6] , \ram[103][5] , \ram[103][4] ,
         \ram[103][3] , \ram[103][2] , \ram[103][1] , \ram[103][0] ,
         \ram[104][7] , \ram[104][6] , \ram[104][5] , \ram[104][4] ,
         \ram[104][3] , \ram[104][2] , \ram[104][1] , \ram[104][0] ,
         \ram[105][7] , \ram[105][6] , \ram[105][5] , \ram[105][4] ,
         \ram[105][3] , \ram[105][2] , \ram[105][1] , \ram[105][0] ,
         \ram[106][7] , \ram[106][6] , \ram[106][5] , \ram[106][4] ,
         \ram[106][3] , \ram[106][2] , \ram[106][1] , \ram[106][0] ,
         \ram[107][7] , \ram[107][6] , \ram[107][5] , \ram[107][4] ,
         \ram[107][3] , \ram[107][2] , \ram[107][1] , \ram[107][0] ,
         \ram[108][7] , \ram[108][6] , \ram[108][5] , \ram[108][4] ,
         \ram[108][3] , \ram[108][2] , \ram[108][1] , \ram[108][0] ,
         \ram[109][7] , \ram[109][6] , \ram[109][5] , \ram[109][4] ,
         \ram[109][3] , \ram[109][2] , \ram[109][1] , \ram[109][0] ,
         \ram[110][7] , \ram[110][6] , \ram[110][5] , \ram[110][4] ,
         \ram[110][3] , \ram[110][2] , \ram[110][1] , \ram[110][0] ,
         \ram[111][7] , \ram[111][6] , \ram[111][5] , \ram[111][4] ,
         \ram[111][3] , \ram[111][2] , \ram[111][1] , \ram[111][0] ,
         \ram[112][7] , \ram[112][6] , \ram[112][5] , \ram[112][4] ,
         \ram[112][3] , \ram[112][2] , \ram[112][1] , \ram[112][0] ,
         \ram[113][7] , \ram[113][6] , \ram[113][5] , \ram[113][4] ,
         \ram[113][3] , \ram[113][2] , \ram[113][1] , \ram[113][0] ,
         \ram[114][7] , \ram[114][6] , \ram[114][5] , \ram[114][4] ,
         \ram[114][3] , \ram[114][2] , \ram[114][1] , \ram[114][0] ,
         \ram[115][7] , \ram[115][6] , \ram[115][5] , \ram[115][4] ,
         \ram[115][3] , \ram[115][2] , \ram[115][1] , \ram[115][0] ,
         \ram[116][7] , \ram[116][6] , \ram[116][5] , \ram[116][4] ,
         \ram[116][3] , \ram[116][2] , \ram[116][1] , \ram[116][0] ,
         \ram[117][7] , \ram[117][6] , \ram[117][5] , \ram[117][4] ,
         \ram[117][3] , \ram[117][2] , \ram[117][1] , \ram[117][0] ,
         \ram[118][7] , \ram[118][6] , \ram[118][5] , \ram[118][4] ,
         \ram[118][3] , \ram[118][2] , \ram[118][1] , \ram[118][0] ,
         \ram[119][7] , \ram[119][6] , \ram[119][5] , \ram[119][4] ,
         \ram[119][3] , \ram[119][2] , \ram[119][1] , \ram[119][0] ,
         \ram[120][7] , \ram[120][6] , \ram[120][5] , \ram[120][4] ,
         \ram[120][3] , \ram[120][2] , \ram[120][1] , \ram[120][0] ,
         \ram[121][7] , \ram[121][6] , \ram[121][5] , \ram[121][4] ,
         \ram[121][3] , \ram[121][2] , \ram[121][1] , \ram[121][0] ,
         \ram[122][7] , \ram[122][6] , \ram[122][5] , \ram[122][4] ,
         \ram[122][3] , \ram[122][2] , \ram[122][1] , \ram[122][0] ,
         \ram[123][7] , \ram[123][6] , \ram[123][5] , \ram[123][4] ,
         \ram[123][3] , \ram[123][2] , \ram[123][1] , \ram[123][0] ,
         \ram[124][7] , \ram[124][6] , \ram[124][5] , \ram[124][4] ,
         \ram[124][3] , \ram[124][2] , \ram[124][1] , \ram[124][0] ,
         \ram[125][7] , \ram[125][6] , \ram[125][5] , \ram[125][4] ,
         \ram[125][3] , \ram[125][2] , \ram[125][1] , \ram[125][0] ,
         \ram[126][7] , \ram[126][6] , \ram[126][5] , \ram[126][4] ,
         \ram[126][3] , \ram[126][2] , \ram[126][1] , \ram[126][0] ,
         \ram[127][7] , \ram[127][6] , \ram[127][5] , \ram[127][4] ,
         \ram[127][3] , \ram[127][2] , \ram[127][1] , \ram[127][0] ,
         \ram[128][7] , \ram[128][6] , \ram[128][5] , \ram[128][4] ,
         \ram[128][3] , \ram[128][2] , \ram[128][1] , \ram[128][0] ,
         \ram[129][7] , \ram[129][6] , \ram[129][5] , \ram[129][4] ,
         \ram[129][3] , \ram[129][2] , \ram[129][1] , \ram[129][0] ,
         \ram[130][7] , \ram[130][6] , \ram[130][5] , \ram[130][4] ,
         \ram[130][3] , \ram[130][2] , \ram[130][1] , \ram[130][0] ,
         \ram[131][7] , \ram[131][6] , \ram[131][5] , \ram[131][4] ,
         \ram[131][3] , \ram[131][2] , \ram[131][1] , \ram[131][0] ,
         \ram[132][7] , \ram[132][6] , \ram[132][5] , \ram[132][4] ,
         \ram[132][3] , \ram[132][2] , \ram[132][1] , \ram[132][0] ,
         \ram[133][7] , \ram[133][6] , \ram[133][5] , \ram[133][4] ,
         \ram[133][3] , \ram[133][2] , \ram[133][1] , \ram[133][0] ,
         \ram[134][7] , \ram[134][6] , \ram[134][5] , \ram[134][4] ,
         \ram[134][3] , \ram[134][2] , \ram[134][1] , \ram[134][0] ,
         \ram[135][7] , \ram[135][6] , \ram[135][5] , \ram[135][4] ,
         \ram[135][3] , \ram[135][2] , \ram[135][1] , \ram[135][0] ,
         \ram[136][7] , \ram[136][6] , \ram[136][5] , \ram[136][4] ,
         \ram[136][3] , \ram[136][2] , \ram[136][1] , \ram[136][0] ,
         \ram[137][7] , \ram[137][6] , \ram[137][5] , \ram[137][4] ,
         \ram[137][3] , \ram[137][2] , \ram[137][1] , \ram[137][0] ,
         \ram[138][7] , \ram[138][6] , \ram[138][5] , \ram[138][4] ,
         \ram[138][3] , \ram[138][2] , \ram[138][1] , \ram[138][0] ,
         \ram[139][7] , \ram[139][6] , \ram[139][5] , \ram[139][4] ,
         \ram[139][3] , \ram[139][2] , \ram[139][1] , \ram[139][0] ,
         \ram[140][7] , \ram[140][6] , \ram[140][5] , \ram[140][4] ,
         \ram[140][3] , \ram[140][2] , \ram[140][1] , \ram[140][0] ,
         \ram[141][7] , \ram[141][6] , \ram[141][5] , \ram[141][4] ,
         \ram[141][3] , \ram[141][2] , \ram[141][1] , \ram[141][0] ,
         \ram[142][7] , \ram[142][6] , \ram[142][5] , \ram[142][4] ,
         \ram[142][3] , \ram[142][2] , \ram[142][1] , \ram[142][0] ,
         \ram[143][7] , \ram[143][6] , \ram[143][5] , \ram[143][4] ,
         \ram[143][3] , \ram[143][2] , \ram[143][1] , \ram[143][0] ,
         \ram[144][7] , \ram[144][6] , \ram[144][5] , \ram[144][4] ,
         \ram[144][3] , \ram[144][2] , \ram[144][1] , \ram[144][0] ,
         \ram[145][7] , \ram[145][6] , \ram[145][5] , \ram[145][4] ,
         \ram[145][3] , \ram[145][2] , \ram[145][1] , \ram[145][0] ,
         \ram[146][7] , \ram[146][6] , \ram[146][5] , \ram[146][4] ,
         \ram[146][3] , \ram[146][2] , \ram[146][1] , \ram[146][0] ,
         \ram[147][7] , \ram[147][6] , \ram[147][5] , \ram[147][4] ,
         \ram[147][3] , \ram[147][2] , \ram[147][1] , \ram[147][0] ,
         \ram[148][7] , \ram[148][6] , \ram[148][5] , \ram[148][4] ,
         \ram[148][3] , \ram[148][2] , \ram[148][1] , \ram[148][0] ,
         \ram[149][7] , \ram[149][6] , \ram[149][5] , \ram[149][4] ,
         \ram[149][3] , \ram[149][2] , \ram[149][1] , \ram[149][0] ,
         \ram[150][7] , \ram[150][6] , \ram[150][5] , \ram[150][4] ,
         \ram[150][3] , \ram[150][2] , \ram[150][1] , \ram[150][0] ,
         \ram[151][7] , \ram[151][6] , \ram[151][5] , \ram[151][4] ,
         \ram[151][3] , \ram[151][2] , \ram[151][1] , \ram[151][0] ,
         \ram[152][7] , \ram[152][6] , \ram[152][5] , \ram[152][4] ,
         \ram[152][3] , \ram[152][2] , \ram[152][1] , \ram[152][0] ,
         \ram[153][7] , \ram[153][6] , \ram[153][5] , \ram[153][4] ,
         \ram[153][3] , \ram[153][2] , \ram[153][1] , \ram[153][0] ,
         \ram[154][7] , \ram[154][6] , \ram[154][5] , \ram[154][4] ,
         \ram[154][3] , \ram[154][2] , \ram[154][1] , \ram[154][0] ,
         \ram[155][7] , \ram[155][6] , \ram[155][5] , \ram[155][4] ,
         \ram[155][3] , \ram[155][2] , \ram[155][1] , \ram[155][0] ,
         \ram[156][7] , \ram[156][6] , \ram[156][5] , \ram[156][4] ,
         \ram[156][3] , \ram[156][2] , \ram[156][1] , \ram[156][0] ,
         \ram[157][7] , \ram[157][6] , \ram[157][5] , \ram[157][4] ,
         \ram[157][3] , \ram[157][2] , \ram[157][1] , \ram[157][0] ,
         \ram[158][7] , \ram[158][6] , \ram[158][5] , \ram[158][4] ,
         \ram[158][3] , \ram[158][2] , \ram[158][1] , \ram[158][0] ,
         \ram[159][7] , \ram[159][6] , \ram[159][5] , \ram[159][4] ,
         \ram[159][3] , \ram[159][2] , \ram[159][1] , \ram[159][0] ,
         \ram[160][7] , \ram[160][6] , \ram[160][5] , \ram[160][4] ,
         \ram[160][3] , \ram[160][2] , \ram[160][1] , \ram[160][0] ,
         \ram[161][7] , \ram[161][6] , \ram[161][5] , \ram[161][4] ,
         \ram[161][3] , \ram[161][2] , \ram[161][1] , \ram[161][0] ,
         \ram[162][7] , \ram[162][6] , \ram[162][5] , \ram[162][4] ,
         \ram[162][3] , \ram[162][2] , \ram[162][1] , \ram[162][0] ,
         \ram[163][7] , \ram[163][6] , \ram[163][5] , \ram[163][4] ,
         \ram[163][3] , \ram[163][2] , \ram[163][1] , \ram[163][0] ,
         \ram[164][7] , \ram[164][6] , \ram[164][5] , \ram[164][4] ,
         \ram[164][3] , \ram[164][2] , \ram[164][1] , \ram[164][0] ,
         \ram[165][7] , \ram[165][6] , \ram[165][5] , \ram[165][4] ,
         \ram[165][3] , \ram[165][2] , \ram[165][1] , \ram[165][0] ,
         \ram[166][7] , \ram[166][6] , \ram[166][5] , \ram[166][4] ,
         \ram[166][3] , \ram[166][2] , \ram[166][1] , \ram[166][0] ,
         \ram[167][7] , \ram[167][6] , \ram[167][5] , \ram[167][4] ,
         \ram[167][3] , \ram[167][2] , \ram[167][1] , \ram[167][0] ,
         \ram[168][7] , \ram[168][6] , \ram[168][5] , \ram[168][4] ,
         \ram[168][3] , \ram[168][2] , \ram[168][1] , \ram[168][0] ,
         \ram[169][7] , \ram[169][6] , \ram[169][5] , \ram[169][4] ,
         \ram[169][3] , \ram[169][2] , \ram[169][1] , \ram[169][0] ,
         \ram[170][7] , \ram[170][6] , \ram[170][5] , \ram[170][4] ,
         \ram[170][3] , \ram[170][2] , \ram[170][1] , \ram[170][0] ,
         \ram[171][7] , \ram[171][6] , \ram[171][5] , \ram[171][4] ,
         \ram[171][3] , \ram[171][2] , \ram[171][1] , \ram[171][0] ,
         \ram[172][7] , \ram[172][6] , \ram[172][5] , \ram[172][4] ,
         \ram[172][3] , \ram[172][2] , \ram[172][1] , \ram[172][0] ,
         \ram[173][7] , \ram[173][6] , \ram[173][5] , \ram[173][4] ,
         \ram[173][3] , \ram[173][2] , \ram[173][1] , \ram[173][0] ,
         \ram[174][7] , \ram[174][6] , \ram[174][5] , \ram[174][4] ,
         \ram[174][3] , \ram[174][2] , \ram[174][1] , \ram[174][0] ,
         \ram[175][7] , \ram[175][6] , \ram[175][5] , \ram[175][4] ,
         \ram[175][3] , \ram[175][2] , \ram[175][1] , \ram[175][0] ,
         \ram[176][7] , \ram[176][6] , \ram[176][5] , \ram[176][4] ,
         \ram[176][3] , \ram[176][2] , \ram[176][1] , \ram[176][0] ,
         \ram[177][7] , \ram[177][6] , \ram[177][5] , \ram[177][4] ,
         \ram[177][3] , \ram[177][2] , \ram[177][1] , \ram[177][0] ,
         \ram[178][7] , \ram[178][6] , \ram[178][5] , \ram[178][4] ,
         \ram[178][3] , \ram[178][2] , \ram[178][1] , \ram[178][0] ,
         \ram[179][7] , \ram[179][6] , \ram[179][5] , \ram[179][4] ,
         \ram[179][3] , \ram[179][2] , \ram[179][1] , \ram[179][0] ,
         \ram[180][7] , \ram[180][6] , \ram[180][5] , \ram[180][4] ,
         \ram[180][3] , \ram[180][2] , \ram[180][1] , \ram[180][0] ,
         \ram[181][7] , \ram[181][6] , \ram[181][5] , \ram[181][4] ,
         \ram[181][3] , \ram[181][2] , \ram[181][1] , \ram[181][0] ,
         \ram[182][7] , \ram[182][6] , \ram[182][5] , \ram[182][4] ,
         \ram[182][3] , \ram[182][2] , \ram[182][1] , \ram[182][0] ,
         \ram[183][7] , \ram[183][6] , \ram[183][5] , \ram[183][4] ,
         \ram[183][3] , \ram[183][2] , \ram[183][1] , \ram[183][0] ,
         \ram[184][7] , \ram[184][6] , \ram[184][5] , \ram[184][4] ,
         \ram[184][3] , \ram[184][2] , \ram[184][1] , \ram[184][0] ,
         \ram[185][7] , \ram[185][6] , \ram[185][5] , \ram[185][4] ,
         \ram[185][3] , \ram[185][2] , \ram[185][1] , \ram[185][0] ,
         \ram[186][7] , \ram[186][6] , \ram[186][5] , \ram[186][4] ,
         \ram[186][3] , \ram[186][2] , \ram[186][1] , \ram[186][0] ,
         \ram[187][7] , \ram[187][6] , \ram[187][5] , \ram[187][4] ,
         \ram[187][3] , \ram[187][2] , \ram[187][1] , \ram[187][0] ,
         \ram[188][7] , \ram[188][6] , \ram[188][5] , \ram[188][4] ,
         \ram[188][3] , \ram[188][2] , \ram[188][1] , \ram[188][0] ,
         \ram[189][7] , \ram[189][6] , \ram[189][5] , \ram[189][4] ,
         \ram[189][3] , \ram[189][2] , \ram[189][1] , \ram[189][0] ,
         \ram[190][7] , \ram[190][6] , \ram[190][5] , \ram[190][4] ,
         \ram[190][3] , \ram[190][2] , \ram[190][1] , \ram[190][0] ,
         \ram[191][7] , \ram[191][6] , \ram[191][5] , \ram[191][4] ,
         \ram[191][3] , \ram[191][2] , \ram[191][1] , \ram[191][0] ,
         \ram[192][7] , \ram[192][6] , \ram[192][5] , \ram[192][4] ,
         \ram[192][3] , \ram[192][2] , \ram[192][1] , \ram[192][0] ,
         \ram[193][7] , \ram[193][6] , \ram[193][5] , \ram[193][4] ,
         \ram[193][3] , \ram[193][2] , \ram[193][1] , \ram[193][0] ,
         \ram[194][7] , \ram[194][6] , \ram[194][5] , \ram[194][4] ,
         \ram[194][3] , \ram[194][2] , \ram[194][1] , \ram[194][0] ,
         \ram[195][7] , \ram[195][6] , \ram[195][5] , \ram[195][4] ,
         \ram[195][3] , \ram[195][2] , \ram[195][1] , \ram[195][0] ,
         \ram[196][7] , \ram[196][6] , \ram[196][5] , \ram[196][4] ,
         \ram[196][3] , \ram[196][2] , \ram[196][1] , \ram[196][0] ,
         \ram[197][7] , \ram[197][6] , \ram[197][5] , \ram[197][4] ,
         \ram[197][3] , \ram[197][2] , \ram[197][1] , \ram[197][0] ,
         \ram[198][7] , \ram[198][6] , \ram[198][5] , \ram[198][4] ,
         \ram[198][3] , \ram[198][2] , \ram[198][1] , \ram[198][0] ,
         \ram[199][7] , \ram[199][6] , \ram[199][5] , \ram[199][4] ,
         \ram[199][3] , \ram[199][2] , \ram[199][1] , \ram[199][0] ,
         \ram[200][7] , \ram[200][6] , \ram[200][5] , \ram[200][4] ,
         \ram[200][3] , \ram[200][2] , \ram[200][1] , \ram[200][0] ,
         \ram[201][7] , \ram[201][6] , \ram[201][5] , \ram[201][4] ,
         \ram[201][3] , \ram[201][2] , \ram[201][1] , \ram[201][0] ,
         \ram[202][7] , \ram[202][6] , \ram[202][5] , \ram[202][4] ,
         \ram[202][3] , \ram[202][2] , \ram[202][1] , \ram[202][0] ,
         \ram[203][7] , \ram[203][6] , \ram[203][5] , \ram[203][4] ,
         \ram[203][3] , \ram[203][2] , \ram[203][1] , \ram[203][0] ,
         \ram[204][7] , \ram[204][6] , \ram[204][5] , \ram[204][4] ,
         \ram[204][3] , \ram[204][2] , \ram[204][1] , \ram[204][0] ,
         \ram[205][7] , \ram[205][6] , \ram[205][5] , \ram[205][4] ,
         \ram[205][3] , \ram[205][2] , \ram[205][1] , \ram[205][0] ,
         \ram[206][7] , \ram[206][6] , \ram[206][5] , \ram[206][4] ,
         \ram[206][3] , \ram[206][2] , \ram[206][1] , \ram[206][0] ,
         \ram[207][7] , \ram[207][6] , \ram[207][5] , \ram[207][4] ,
         \ram[207][3] , \ram[207][2] , \ram[207][1] , \ram[207][0] ,
         \ram[208][7] , \ram[208][6] , \ram[208][5] , \ram[208][4] ,
         \ram[208][3] , \ram[208][2] , \ram[208][1] , \ram[208][0] ,
         \ram[209][7] , \ram[209][6] , \ram[209][5] , \ram[209][4] ,
         \ram[209][3] , \ram[209][2] , \ram[209][1] , \ram[209][0] ,
         \ram[210][7] , \ram[210][6] , \ram[210][5] , \ram[210][4] ,
         \ram[210][3] , \ram[210][2] , \ram[210][1] , \ram[210][0] ,
         \ram[211][7] , \ram[211][6] , \ram[211][5] , \ram[211][4] ,
         \ram[211][3] , \ram[211][2] , \ram[211][1] , \ram[211][0] ,
         \ram[212][7] , \ram[212][6] , \ram[212][5] , \ram[212][4] ,
         \ram[212][3] , \ram[212][2] , \ram[212][1] , \ram[212][0] ,
         \ram[213][7] , \ram[213][6] , \ram[213][5] , \ram[213][4] ,
         \ram[213][3] , \ram[213][2] , \ram[213][1] , \ram[213][0] ,
         \ram[214][7] , \ram[214][6] , \ram[214][5] , \ram[214][4] ,
         \ram[214][3] , \ram[214][2] , \ram[214][1] , \ram[214][0] ,
         \ram[215][7] , \ram[215][6] , \ram[215][5] , \ram[215][4] ,
         \ram[215][3] , \ram[215][2] , \ram[215][1] , \ram[215][0] ,
         \ram[216][7] , \ram[216][6] , \ram[216][5] , \ram[216][4] ,
         \ram[216][3] , \ram[216][2] , \ram[216][1] , \ram[216][0] ,
         \ram[217][7] , \ram[217][6] , \ram[217][5] , \ram[217][4] ,
         \ram[217][3] , \ram[217][2] , \ram[217][1] , \ram[217][0] ,
         \ram[218][7] , \ram[218][6] , \ram[218][5] , \ram[218][4] ,
         \ram[218][3] , \ram[218][2] , \ram[218][1] , \ram[218][0] ,
         \ram[219][7] , \ram[219][6] , \ram[219][5] , \ram[219][4] ,
         \ram[219][3] , \ram[219][2] , \ram[219][1] , \ram[219][0] ,
         \ram[220][7] , \ram[220][6] , \ram[220][5] , \ram[220][4] ,
         \ram[220][3] , \ram[220][2] , \ram[220][1] , \ram[220][0] ,
         \ram[221][7] , \ram[221][6] , \ram[221][5] , \ram[221][4] ,
         \ram[221][3] , \ram[221][2] , \ram[221][1] , \ram[221][0] ,
         \ram[222][7] , \ram[222][6] , \ram[222][5] , \ram[222][4] ,
         \ram[222][3] , \ram[222][2] , \ram[222][1] , \ram[222][0] ,
         \ram[223][7] , \ram[223][6] , \ram[223][5] , \ram[223][4] ,
         \ram[223][3] , \ram[223][2] , \ram[223][1] , \ram[223][0] ,
         \ram[224][7] , \ram[224][6] , \ram[224][5] , \ram[224][4] ,
         \ram[224][3] , \ram[224][2] , \ram[224][1] , \ram[224][0] ,
         \ram[225][7] , \ram[225][6] , \ram[225][5] , \ram[225][4] ,
         \ram[225][3] , \ram[225][2] , \ram[225][1] , \ram[225][0] ,
         \ram[226][7] , \ram[226][6] , \ram[226][5] , \ram[226][4] ,
         \ram[226][3] , \ram[226][2] , \ram[226][1] , \ram[226][0] ,
         \ram[227][7] , \ram[227][6] , \ram[227][5] , \ram[227][4] ,
         \ram[227][3] , \ram[227][2] , \ram[227][1] , \ram[227][0] ,
         \ram[228][7] , \ram[228][6] , \ram[228][5] , \ram[228][4] ,
         \ram[228][3] , \ram[228][2] , \ram[228][1] , \ram[228][0] ,
         \ram[229][7] , \ram[229][6] , \ram[229][5] , \ram[229][4] ,
         \ram[229][3] , \ram[229][2] , \ram[229][1] , \ram[229][0] ,
         \ram[230][7] , \ram[230][6] , \ram[230][5] , \ram[230][4] ,
         \ram[230][3] , \ram[230][2] , \ram[230][1] , \ram[230][0] ,
         \ram[231][7] , \ram[231][6] , \ram[231][5] , \ram[231][4] ,
         \ram[231][3] , \ram[231][2] , \ram[231][1] , \ram[231][0] ,
         \ram[232][7] , \ram[232][6] , \ram[232][5] , \ram[232][4] ,
         \ram[232][3] , \ram[232][2] , \ram[232][1] , \ram[232][0] ,
         \ram[233][7] , \ram[233][6] , \ram[233][5] , \ram[233][4] ,
         \ram[233][3] , \ram[233][2] , \ram[233][1] , \ram[233][0] ,
         \ram[234][7] , \ram[234][6] , \ram[234][5] , \ram[234][4] ,
         \ram[234][3] , \ram[234][2] , \ram[234][1] , \ram[234][0] ,
         \ram[235][7] , \ram[235][6] , \ram[235][5] , \ram[235][4] ,
         \ram[235][3] , \ram[235][2] , \ram[235][1] , \ram[235][0] ,
         \ram[236][7] , \ram[236][6] , \ram[236][5] , \ram[236][4] ,
         \ram[236][3] , \ram[236][2] , \ram[236][1] , \ram[236][0] ,
         \ram[237][7] , \ram[237][6] , \ram[237][5] , \ram[237][4] ,
         \ram[237][3] , \ram[237][2] , \ram[237][1] , \ram[237][0] ,
         \ram[238][7] , \ram[238][6] , \ram[238][5] , \ram[238][4] ,
         \ram[238][3] , \ram[238][2] , \ram[238][1] , \ram[238][0] ,
         \ram[239][7] , \ram[239][6] , \ram[239][5] , \ram[239][4] ,
         \ram[239][3] , \ram[239][2] , \ram[239][1] , \ram[239][0] ,
         \ram[240][7] , \ram[240][6] , \ram[240][5] , \ram[240][4] ,
         \ram[240][3] , \ram[240][2] , \ram[240][1] , \ram[240][0] ,
         \ram[241][7] , \ram[241][6] , \ram[241][5] , \ram[241][4] ,
         \ram[241][3] , \ram[241][2] , \ram[241][1] , \ram[241][0] ,
         \ram[242][7] , \ram[242][6] , \ram[242][5] , \ram[242][4] ,
         \ram[242][3] , \ram[242][2] , \ram[242][1] , \ram[242][0] ,
         \ram[243][7] , \ram[243][6] , \ram[243][5] , \ram[243][4] ,
         \ram[243][3] , \ram[243][2] , \ram[243][1] , \ram[243][0] ,
         \ram[244][7] , \ram[244][6] , \ram[244][5] , \ram[244][4] ,
         \ram[244][3] , \ram[244][2] , \ram[244][1] , \ram[244][0] ,
         \ram[245][7] , \ram[245][6] , \ram[245][5] , \ram[245][4] ,
         \ram[245][3] , \ram[245][2] , \ram[245][1] , \ram[245][0] ,
         \ram[246][7] , \ram[246][6] , \ram[246][5] , \ram[246][4] ,
         \ram[246][3] , \ram[246][2] , \ram[246][1] , \ram[246][0] ,
         \ram[247][7] , \ram[247][6] , \ram[247][5] , \ram[247][4] ,
         \ram[247][3] , \ram[247][2] , \ram[247][1] , \ram[247][0] ,
         \ram[248][7] , \ram[248][6] , \ram[248][5] , \ram[248][4] ,
         \ram[248][3] , \ram[248][2] , \ram[248][1] , \ram[248][0] ,
         \ram[249][7] , \ram[249][6] , \ram[249][5] , \ram[249][4] ,
         \ram[249][3] , \ram[249][2] , \ram[249][1] , \ram[249][0] ,
         \ram[250][7] , \ram[250][6] , \ram[250][5] , \ram[250][4] ,
         \ram[250][3] , \ram[250][2] , \ram[250][1] , \ram[250][0] ,
         \ram[251][7] , \ram[251][6] , \ram[251][5] , \ram[251][4] ,
         \ram[251][3] , \ram[251][2] , \ram[251][1] , \ram[251][0] ,
         \ram[252][7] , \ram[252][6] , \ram[252][5] , \ram[252][4] ,
         \ram[252][3] , \ram[252][2] , \ram[252][1] , \ram[252][0] ,
         \ram[253][7] , \ram[253][6] , \ram[253][5] , \ram[253][4] ,
         \ram[253][3] , \ram[253][2] , \ram[253][1] , \ram[253][0] ,
         \ram[254][7] , \ram[254][6] , \ram[254][5] , \ram[254][4] ,
         \ram[254][3] , \ram[254][2] , \ram[254][1] , \ram[254][0] ,
         \ram[255][7] , \ram[255][6] , \ram[255][5] , \ram[255][4] ,
         \ram[255][3] , \ram[255][2] , \ram[255][1] , \ram[255][0] , n1, n3,
         n4, n5, n7, n8, n10, n11, n13, n14, n16, n17, n19, n20, n22, n23, n25,
         n26, n28, n29, n31, n32, n34, n35, n37, n38, n40, n41, n43, n44, n46,
         n47, n49, n50, n52, n53, n55, n56, n58, n59, n61, n62, n64, n65, n67,
         n68, n70, n71, n73, n74, n76, n77, n79, n80, n82, n83, n85, n86, n88,
         n89, n91, n92, n94, n95, n97, n98, n100, n101, n103, n104, n106, n107,
         n109, n110, n112, n113, n115, n116, n118, n119, n121, n122, n124,
         n125, n127, n128, n130, n131, n133, n134, n136, n137, n139, n140,
         n142, n143, n145, n146, n148, n149, n151, n152, n154, n155, n157,
         n158, n160, n161, n163, n164, n166, n167, n169, n170, n172, n173,
         n175, n176, n178, n179, n181, n182, n184, n185, n187, n188, n190,
         n191, n193, n194, n196, n197, n199, n200, n202, n203, n205, n206,
         n208, n209, n211, n212, n214, n215, n217, n218, n220, n221, n223,
         n224, n226, n227, n229, n230, n232, n233, n235, n236, n238, n239,
         n241, n242, n244, n245, n247, n248, n250, n251, n253, n254, n256,
         n257, n259, n260, n262, n263, n265, n266, n268, n269, n271, n272,
         n274, n275, n277, n278, n280, n281, n283, n284, n286, n287, n289,
         n290, n292, n293, n295, n296, n298, n299, n301, n302, n304, n305,
         n307, n308, n310, n311, n313, n314, n316, n317, n319, n320, n322,
         n323, n325, n326, n328, n329, n331, n332, n334, n335, n337, n338,
         n340, n341, n343, n344, n346, n347, n349, n350, n352, n353, n355,
         n356, n358, n359, n361, n362, n364, n365, n367, n368, n370, n371,
         n373, n374, n376, n377, n379, n380, n382, n383, n385, n386, n388,
         n389, n391, n392, n394, n395, n397, n398, n400, n401, n403, n404,
         n406, n407, n409, n410, n412, n413, n415, n416, n418, n419, n421,
         n422, n424, n425, n427, n428, n430, n431, n433, n434, n436, n437,
         n439, n440, n442, n443, n445, n446, n448, n449, n451, n452, n454,
         n455, n457, n458, n460, n461, n463, n464, n466, n467, n469, n470,
         n472, n473, n475, n476, n478, n479, n481, n482, n484, n485, n487,
         n488, n490, n491, n493, n494, n496, n497, n499, n500, n502, n503,
         n505, n506, n508, n509, n511, n512, n514, n515, n517, n518, n520,
         n521, n523, n524, n526, n527, n529, n530, n532, n533, n535, n536,
         n538, n539, n541, n542, n544, n545, n547, n548, n550, n551, n553,
         n554, n556, n557, n559, n560, n562, n563, n565, n566, n568, n569,
         n571, n572, n574, n575, n577, n578, n580, n581, n583, n584, n586,
         n587, n589, n590, n592, n593, n595, n596, n598, n599, n601, n602,
         n604, n605, n607, n608, n610, n611, n613, n614, n616, n617, n619,
         n620, n622, n623, n625, n626, n628, n629, n631, n632, n634, n635,
         n637, n638, n640, n641, n643, n644, n646, n647, n649, n650, n652,
         n653, n655, n656, n658, n659, n661, n662, n664, n665, n667, n668,
         n670, n671, n673, n674, n676, n677, n679, n680, n682, n683, n685,
         n686, n688, n689, n691, n692, n694, n695, n697, n698, n700, n701,
         n703, n704, n706, n707, n709, n710, n712, n713, n715, n716, n718,
         n719, n721, n722, n724, n725, n727, n728, n730, n731, n733, n734,
         n736, n737, n739, n740, n742, n743, n745, n746, n748, n749, n751,
         n752, n754, n755, n757, n758, n760, n761, n763, n764, n766, n767,
         n769, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2017, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n2, n6, n9, n12, n15,
         n18, n21, n24, n27, n30, n33, n36, n39, n42, n45, n48, n51, n54, n57,
         n60, n63, n66, n69, n72, n75, n78, n81, n84, n87, n90, n93, n96, n99,
         n102, n105, n108, n111, n114, n117, n120, n123, n126, n129, n132,
         n135, n138, n141, n144, n147, n150, n153, n156, n159, n162, n165,
         n168, n171, n174, n177, n180, n183, n186, n189, n192, n195, n198,
         n201, n204, n207, n210, n213, n216, n219, n222, n225, n228, n231,
         n234, n237, n240, n243, n246, n249, n252, n255, n258, n261, n264,
         n267, n270, n273, n276, n279, n282, n285, n288, n291, n294, n297,
         n300, n303, n306, n309, n312, n315, n318, n321, n324, n327, n330,
         n333, n336, n339, n342, n345, n348, n351, n354, n357, n360, n363,
         n366, n369, n372, n375, n378, n381, n384, n387, n390, n393, n396,
         n399, n402, n405, n408, n411, n414, n417, n420, n423, n426, n429,
         n432, n435, n438, n441, n444, n447, n450, n453, n456, n459, n462,
         n465, n468, n471, n474, n477, n480, n483, n486, n489, n492, n495,
         n498, n501, n504, n507, n510, n513, n516, n519, n522, n525, n528,
         n531, n534, n537, n540, n543, n546, n549, n552, n555, n558, n561,
         n564, n567, n570, n573, n576, n579, n582, n585, n588, n591, n594,
         n597, n600, n603, n606, n609, n612, n615, n618, n621, n624, n627,
         n630, n633, n636, n639, n642, n645, n648, n651, n654, n657, n660,
         n663, n666, n669, n672, n675, n678, n681, n684, n687, n690, n693,
         n696, n699, n702, n705, n708, n711, n714, n717, n720, n723, n726,
         n729, n732, n735, n738, n741, n744, n747, n750, n753, n756, n759,
         n762, n765, n768, n770, n1974, n1975, n2006, n2007, n2015, n2016,
         n2018, n2019, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175;

  DFFNX1 \ram_reg[0][7]  ( .D(n4075), .CLK(clk), .Q(\ram[0][7] ) );
  DFFNX1 \ram_reg[0][6]  ( .D(n4074), .CLK(clk), .Q(\ram[0][6] ) );
  DFFNX1 \ram_reg[0][5]  ( .D(n4073), .CLK(clk), .Q(\ram[0][5] ) );
  DFFNX1 \ram_reg[0][4]  ( .D(n4072), .CLK(clk), .Q(\ram[0][4] ) );
  DFFNX1 \ram_reg[0][3]  ( .D(n4071), .CLK(clk), .Q(\ram[0][3] ) );
  DFFNX1 \ram_reg[0][2]  ( .D(n4070), .CLK(clk), .Q(\ram[0][2] ) );
  DFFNX1 \ram_reg[0][1]  ( .D(n4069), .CLK(clk), .Q(\ram[0][1] ) );
  DFFNX1 \ram_reg[0][0]  ( .D(n4068), .CLK(clk), .Q(\ram[0][0] ) );
  DFFNX1 \ram_reg[1][7]  ( .D(n4067), .CLK(clk), .Q(\ram[1][7] ) );
  DFFNX1 \ram_reg[1][6]  ( .D(n4066), .CLK(clk), .Q(\ram[1][6] ) );
  DFFNX1 \ram_reg[1][5]  ( .D(n4065), .CLK(clk), .Q(\ram[1][5] ) );
  DFFNX1 \ram_reg[1][4]  ( .D(n4064), .CLK(clk), .Q(\ram[1][4] ) );
  DFFNX1 \ram_reg[1][3]  ( .D(n4063), .CLK(clk), .Q(\ram[1][3] ) );
  DFFNX1 \ram_reg[1][2]  ( .D(n4062), .CLK(clk), .Q(\ram[1][2] ) );
  DFFNX1 \ram_reg[1][1]  ( .D(n4061), .CLK(clk), .Q(\ram[1][1] ) );
  DFFNX1 \ram_reg[1][0]  ( .D(n4060), .CLK(clk), .Q(\ram[1][0] ) );
  DFFNX1 \ram_reg[2][7]  ( .D(n4059), .CLK(clk), .Q(\ram[2][7] ) );
  DFFNX1 \ram_reg[2][6]  ( .D(n4058), .CLK(clk), .Q(\ram[2][6] ) );
  DFFNX1 \ram_reg[2][5]  ( .D(n4057), .CLK(clk), .Q(\ram[2][5] ) );
  DFFNX1 \ram_reg[2][4]  ( .D(n4056), .CLK(clk), .Q(\ram[2][4] ) );
  DFFNX1 \ram_reg[2][3]  ( .D(n4055), .CLK(clk), .Q(\ram[2][3] ) );
  DFFNX1 \ram_reg[2][2]  ( .D(n4054), .CLK(clk), .Q(\ram[2][2] ) );
  DFFNX1 \ram_reg[2][1]  ( .D(n4053), .CLK(clk), .Q(\ram[2][1] ) );
  DFFNX1 \ram_reg[2][0]  ( .D(n4052), .CLK(clk), .Q(\ram[2][0] ) );
  DFFNX1 \ram_reg[3][7]  ( .D(n4051), .CLK(clk), .Q(\ram[3][7] ) );
  DFFNX1 \ram_reg[3][6]  ( .D(n4050), .CLK(clk), .Q(\ram[3][6] ) );
  DFFNX1 \ram_reg[3][5]  ( .D(n4049), .CLK(clk), .Q(\ram[3][5] ) );
  DFFNX1 \ram_reg[3][4]  ( .D(n4048), .CLK(clk), .Q(\ram[3][4] ) );
  DFFNX1 \ram_reg[3][3]  ( .D(n4047), .CLK(clk), .Q(\ram[3][3] ) );
  DFFNX1 \ram_reg[3][2]  ( .D(n4046), .CLK(clk), .Q(\ram[3][2] ) );
  DFFNX1 \ram_reg[3][1]  ( .D(n4045), .CLK(clk), .Q(\ram[3][1] ) );
  DFFNX1 \ram_reg[3][0]  ( .D(n4044), .CLK(clk), .Q(\ram[3][0] ) );
  DFFNX1 \ram_reg[4][7]  ( .D(n4043), .CLK(clk), .Q(\ram[4][7] ) );
  DFFNX1 \ram_reg[4][6]  ( .D(n4042), .CLK(clk), .Q(\ram[4][6] ) );
  DFFNX1 \ram_reg[4][5]  ( .D(n4041), .CLK(clk), .Q(\ram[4][5] ) );
  DFFNX1 \ram_reg[4][4]  ( .D(n4040), .CLK(clk), .Q(\ram[4][4] ) );
  DFFNX1 \ram_reg[4][3]  ( .D(n4039), .CLK(clk), .Q(\ram[4][3] ) );
  DFFNX1 \ram_reg[4][2]  ( .D(n4038), .CLK(clk), .Q(\ram[4][2] ) );
  DFFNX1 \ram_reg[4][1]  ( .D(n4037), .CLK(clk), .Q(\ram[4][1] ) );
  DFFNX1 \ram_reg[4][0]  ( .D(n4036), .CLK(clk), .Q(\ram[4][0] ) );
  DFFNX1 \ram_reg[5][7]  ( .D(n4035), .CLK(clk), .Q(\ram[5][7] ) );
  DFFNX1 \ram_reg[5][6]  ( .D(n4034), .CLK(clk), .Q(\ram[5][6] ) );
  DFFNX1 \ram_reg[5][5]  ( .D(n4033), .CLK(clk), .Q(\ram[5][5] ) );
  DFFNX1 \ram_reg[5][4]  ( .D(n4032), .CLK(clk), .Q(\ram[5][4] ) );
  DFFNX1 \ram_reg[5][3]  ( .D(n4031), .CLK(clk), .Q(\ram[5][3] ) );
  DFFNX1 \ram_reg[5][2]  ( .D(n4030), .CLK(clk), .Q(\ram[5][2] ) );
  DFFNX1 \ram_reg[5][1]  ( .D(n4029), .CLK(clk), .Q(\ram[5][1] ) );
  DFFNX1 \ram_reg[5][0]  ( .D(n4028), .CLK(clk), .Q(\ram[5][0] ) );
  DFFNX1 \ram_reg[6][7]  ( .D(n4027), .CLK(clk), .Q(\ram[6][7] ) );
  DFFNX1 \ram_reg[6][6]  ( .D(n4026), .CLK(clk), .Q(\ram[6][6] ) );
  DFFNX1 \ram_reg[6][5]  ( .D(n4025), .CLK(clk), .Q(\ram[6][5] ) );
  DFFNX1 \ram_reg[6][4]  ( .D(n4024), .CLK(clk), .Q(\ram[6][4] ) );
  DFFNX1 \ram_reg[6][3]  ( .D(n4023), .CLK(clk), .Q(\ram[6][3] ) );
  DFFNX1 \ram_reg[6][2]  ( .D(n4022), .CLK(clk), .Q(\ram[6][2] ) );
  DFFNX1 \ram_reg[6][1]  ( .D(n4021), .CLK(clk), .Q(\ram[6][1] ) );
  DFFNX1 \ram_reg[6][0]  ( .D(n4020), .CLK(clk), .Q(\ram[6][0] ) );
  DFFNX1 \ram_reg[7][7]  ( .D(n4019), .CLK(clk), .Q(\ram[7][7] ) );
  DFFNX1 \ram_reg[7][6]  ( .D(n4018), .CLK(clk), .Q(\ram[7][6] ) );
  DFFNX1 \ram_reg[7][5]  ( .D(n4017), .CLK(clk), .Q(\ram[7][5] ) );
  DFFNX1 \ram_reg[7][4]  ( .D(n4016), .CLK(clk), .Q(\ram[7][4] ) );
  DFFNX1 \ram_reg[7][3]  ( .D(n4015), .CLK(clk), .Q(\ram[7][3] ) );
  DFFNX1 \ram_reg[7][2]  ( .D(n4014), .CLK(clk), .Q(\ram[7][2] ) );
  DFFNX1 \ram_reg[7][1]  ( .D(n4013), .CLK(clk), .Q(\ram[7][1] ) );
  DFFNX1 \ram_reg[7][0]  ( .D(n4012), .CLK(clk), .Q(\ram[7][0] ) );
  DFFNX1 \ram_reg[8][7]  ( .D(n4011), .CLK(clk), .Q(\ram[8][7] ) );
  DFFNX1 \ram_reg[8][6]  ( .D(n4010), .CLK(clk), .Q(\ram[8][6] ) );
  DFFNX1 \ram_reg[8][5]  ( .D(n4009), .CLK(clk), .Q(\ram[8][5] ) );
  DFFNX1 \ram_reg[8][4]  ( .D(n4008), .CLK(clk), .Q(\ram[8][4] ) );
  DFFNX1 \ram_reg[8][3]  ( .D(n4007), .CLK(clk), .Q(\ram[8][3] ) );
  DFFNX1 \ram_reg[8][2]  ( .D(n4006), .CLK(clk), .Q(\ram[8][2] ) );
  DFFNX1 \ram_reg[8][1]  ( .D(n4005), .CLK(clk), .Q(\ram[8][1] ) );
  DFFNX1 \ram_reg[8][0]  ( .D(n4004), .CLK(clk), .Q(\ram[8][0] ) );
  DFFNX1 \ram_reg[9][7]  ( .D(n4003), .CLK(clk), .Q(\ram[9][7] ) );
  DFFNX1 \ram_reg[9][6]  ( .D(n4002), .CLK(clk), .Q(\ram[9][6] ) );
  DFFNX1 \ram_reg[9][5]  ( .D(n4001), .CLK(clk), .Q(\ram[9][5] ) );
  DFFNX1 \ram_reg[9][4]  ( .D(n4000), .CLK(clk), .Q(\ram[9][4] ) );
  DFFNX1 \ram_reg[9][3]  ( .D(n3999), .CLK(clk), .Q(\ram[9][3] ) );
  DFFNX1 \ram_reg[9][2]  ( .D(n3998), .CLK(clk), .Q(\ram[9][2] ) );
  DFFNX1 \ram_reg[9][1]  ( .D(n3997), .CLK(clk), .Q(\ram[9][1] ) );
  DFFNX1 \ram_reg[9][0]  ( .D(n3996), .CLK(clk), .Q(\ram[9][0] ) );
  DFFNX1 \ram_reg[10][7]  ( .D(n3995), .CLK(clk), .Q(\ram[10][7] ) );
  DFFNX1 \ram_reg[10][6]  ( .D(n3994), .CLK(clk), .Q(\ram[10][6] ) );
  DFFNX1 \ram_reg[10][5]  ( .D(n3993), .CLK(clk), .Q(\ram[10][5] ) );
  DFFNX1 \ram_reg[10][4]  ( .D(n3992), .CLK(clk), .Q(\ram[10][4] ) );
  DFFNX1 \ram_reg[10][3]  ( .D(n3991), .CLK(clk), .Q(\ram[10][3] ) );
  DFFNX1 \ram_reg[10][2]  ( .D(n3990), .CLK(clk), .Q(\ram[10][2] ) );
  DFFNX1 \ram_reg[10][1]  ( .D(n3989), .CLK(clk), .Q(\ram[10][1] ) );
  DFFNX1 \ram_reg[10][0]  ( .D(n3988), .CLK(clk), .Q(\ram[10][0] ) );
  DFFNX1 \ram_reg[11][7]  ( .D(n3987), .CLK(clk), .Q(\ram[11][7] ) );
  DFFNX1 \ram_reg[11][6]  ( .D(n3986), .CLK(clk), .Q(\ram[11][6] ) );
  DFFNX1 \ram_reg[11][5]  ( .D(n3985), .CLK(clk), .Q(\ram[11][5] ) );
  DFFNX1 \ram_reg[11][4]  ( .D(n3984), .CLK(clk), .Q(\ram[11][4] ) );
  DFFNX1 \ram_reg[11][3]  ( .D(n3983), .CLK(clk), .Q(\ram[11][3] ) );
  DFFNX1 \ram_reg[11][2]  ( .D(n3982), .CLK(clk), .Q(\ram[11][2] ) );
  DFFNX1 \ram_reg[11][1]  ( .D(n3981), .CLK(clk), .Q(\ram[11][1] ) );
  DFFNX1 \ram_reg[11][0]  ( .D(n3980), .CLK(clk), .Q(\ram[11][0] ) );
  DFFNX1 \ram_reg[12][7]  ( .D(n3979), .CLK(clk), .Q(\ram[12][7] ) );
  DFFNX1 \ram_reg[12][6]  ( .D(n3978), .CLK(clk), .Q(\ram[12][6] ) );
  DFFNX1 \ram_reg[12][5]  ( .D(n3977), .CLK(clk), .Q(\ram[12][5] ) );
  DFFNX1 \ram_reg[12][4]  ( .D(n3976), .CLK(clk), .Q(\ram[12][4] ) );
  DFFNX1 \ram_reg[12][3]  ( .D(n3975), .CLK(clk), .Q(\ram[12][3] ) );
  DFFNX1 \ram_reg[12][2]  ( .D(n3974), .CLK(clk), .Q(\ram[12][2] ) );
  DFFNX1 \ram_reg[12][1]  ( .D(n3973), .CLK(clk), .Q(\ram[12][1] ) );
  DFFNX1 \ram_reg[12][0]  ( .D(n3972), .CLK(clk), .Q(\ram[12][0] ) );
  DFFNX1 \ram_reg[13][7]  ( .D(n3971), .CLK(clk), .Q(\ram[13][7] ) );
  DFFNX1 \ram_reg[13][6]  ( .D(n3970), .CLK(clk), .Q(\ram[13][6] ) );
  DFFNX1 \ram_reg[13][5]  ( .D(n3969), .CLK(clk), .Q(\ram[13][5] ) );
  DFFNX1 \ram_reg[13][4]  ( .D(n3968), .CLK(clk), .Q(\ram[13][4] ) );
  DFFNX1 \ram_reg[13][3]  ( .D(n3967), .CLK(clk), .Q(\ram[13][3] ) );
  DFFNX1 \ram_reg[13][2]  ( .D(n3966), .CLK(clk), .Q(\ram[13][2] ) );
  DFFNX1 \ram_reg[13][1]  ( .D(n3965), .CLK(clk), .Q(\ram[13][1] ) );
  DFFNX1 \ram_reg[13][0]  ( .D(n3964), .CLK(clk), .Q(\ram[13][0] ) );
  DFFNX1 \ram_reg[14][7]  ( .D(n3963), .CLK(clk), .Q(\ram[14][7] ) );
  DFFNX1 \ram_reg[14][6]  ( .D(n3962), .CLK(clk), .Q(\ram[14][6] ) );
  DFFNX1 \ram_reg[14][5]  ( .D(n3961), .CLK(clk), .Q(\ram[14][5] ) );
  DFFNX1 \ram_reg[14][4]  ( .D(n3960), .CLK(clk), .Q(\ram[14][4] ) );
  DFFNX1 \ram_reg[14][3]  ( .D(n3959), .CLK(clk), .Q(\ram[14][3] ) );
  DFFNX1 \ram_reg[14][2]  ( .D(n3958), .CLK(clk), .Q(\ram[14][2] ) );
  DFFNX1 \ram_reg[14][1]  ( .D(n3957), .CLK(clk), .Q(\ram[14][1] ) );
  DFFNX1 \ram_reg[14][0]  ( .D(n3956), .CLK(clk), .Q(\ram[14][0] ) );
  DFFNX1 \ram_reg[15][7]  ( .D(n3955), .CLK(clk), .Q(\ram[15][7] ) );
  DFFNX1 \ram_reg[15][6]  ( .D(n3954), .CLK(clk), .Q(\ram[15][6] ) );
  DFFNX1 \ram_reg[15][5]  ( .D(n3953), .CLK(clk), .Q(\ram[15][5] ) );
  DFFNX1 \ram_reg[15][4]  ( .D(n3952), .CLK(clk), .Q(\ram[15][4] ) );
  DFFNX1 \ram_reg[15][3]  ( .D(n3951), .CLK(clk), .Q(\ram[15][3] ) );
  DFFNX1 \ram_reg[15][2]  ( .D(n3950), .CLK(clk), .Q(\ram[15][2] ) );
  DFFNX1 \ram_reg[15][1]  ( .D(n3949), .CLK(clk), .Q(\ram[15][1] ) );
  DFFNX1 \ram_reg[15][0]  ( .D(n3948), .CLK(clk), .Q(\ram[15][0] ) );
  DFFNX1 \ram_reg[16][7]  ( .D(n3947), .CLK(clk), .Q(\ram[16][7] ) );
  DFFNX1 \ram_reg[16][6]  ( .D(n3946), .CLK(clk), .Q(\ram[16][6] ) );
  DFFNX1 \ram_reg[16][5]  ( .D(n3945), .CLK(clk), .Q(\ram[16][5] ) );
  DFFNX1 \ram_reg[16][4]  ( .D(n3944), .CLK(clk), .Q(\ram[16][4] ) );
  DFFNX1 \ram_reg[16][3]  ( .D(n3943), .CLK(clk), .Q(\ram[16][3] ) );
  DFFNX1 \ram_reg[16][2]  ( .D(n3942), .CLK(clk), .Q(\ram[16][2] ) );
  DFFNX1 \ram_reg[16][1]  ( .D(n3941), .CLK(clk), .Q(\ram[16][1] ) );
  DFFNX1 \ram_reg[16][0]  ( .D(n3940), .CLK(clk), .Q(\ram[16][0] ) );
  DFFNX1 \ram_reg[17][7]  ( .D(n3939), .CLK(clk), .Q(\ram[17][7] ) );
  DFFNX1 \ram_reg[17][6]  ( .D(n3938), .CLK(clk), .Q(\ram[17][6] ) );
  DFFNX1 \ram_reg[17][5]  ( .D(n3937), .CLK(clk), .Q(\ram[17][5] ) );
  DFFNX1 \ram_reg[17][4]  ( .D(n3936), .CLK(clk), .Q(\ram[17][4] ) );
  DFFNX1 \ram_reg[17][3]  ( .D(n3935), .CLK(clk), .Q(\ram[17][3] ) );
  DFFNX1 \ram_reg[17][2]  ( .D(n3934), .CLK(clk), .Q(\ram[17][2] ) );
  DFFNX1 \ram_reg[17][1]  ( .D(n3933), .CLK(clk), .Q(\ram[17][1] ) );
  DFFNX1 \ram_reg[17][0]  ( .D(n3932), .CLK(clk), .Q(\ram[17][0] ) );
  DFFNX1 \ram_reg[18][7]  ( .D(n3931), .CLK(clk), .Q(\ram[18][7] ) );
  DFFNX1 \ram_reg[18][6]  ( .D(n3930), .CLK(clk), .Q(\ram[18][6] ) );
  DFFNX1 \ram_reg[18][5]  ( .D(n3929), .CLK(clk), .Q(\ram[18][5] ) );
  DFFNX1 \ram_reg[18][4]  ( .D(n3928), .CLK(clk), .Q(\ram[18][4] ) );
  DFFNX1 \ram_reg[18][3]  ( .D(n3927), .CLK(clk), .Q(\ram[18][3] ) );
  DFFNX1 \ram_reg[18][2]  ( .D(n3926), .CLK(clk), .Q(\ram[18][2] ) );
  DFFNX1 \ram_reg[18][1]  ( .D(n3925), .CLK(clk), .Q(\ram[18][1] ) );
  DFFNX1 \ram_reg[18][0]  ( .D(n3924), .CLK(clk), .Q(\ram[18][0] ) );
  DFFNX1 \ram_reg[19][7]  ( .D(n3923), .CLK(clk), .Q(\ram[19][7] ) );
  DFFNX1 \ram_reg[19][6]  ( .D(n3922), .CLK(clk), .Q(\ram[19][6] ) );
  DFFNX1 \ram_reg[19][5]  ( .D(n3921), .CLK(clk), .Q(\ram[19][5] ) );
  DFFNX1 \ram_reg[19][4]  ( .D(n3920), .CLK(clk), .Q(\ram[19][4] ) );
  DFFNX1 \ram_reg[19][3]  ( .D(n3919), .CLK(clk), .Q(\ram[19][3] ) );
  DFFNX1 \ram_reg[19][2]  ( .D(n3918), .CLK(clk), .Q(\ram[19][2] ) );
  DFFNX1 \ram_reg[19][1]  ( .D(n3917), .CLK(clk), .Q(\ram[19][1] ) );
  DFFNX1 \ram_reg[19][0]  ( .D(n3916), .CLK(clk), .Q(\ram[19][0] ) );
  DFFNX1 \ram_reg[20][7]  ( .D(n3915), .CLK(clk), .Q(\ram[20][7] ) );
  DFFNX1 \ram_reg[20][6]  ( .D(n3914), .CLK(clk), .Q(\ram[20][6] ) );
  DFFNX1 \ram_reg[20][5]  ( .D(n3913), .CLK(clk), .Q(\ram[20][5] ) );
  DFFNX1 \ram_reg[20][4]  ( .D(n3912), .CLK(clk), .Q(\ram[20][4] ) );
  DFFNX1 \ram_reg[20][3]  ( .D(n3911), .CLK(clk), .Q(\ram[20][3] ) );
  DFFNX1 \ram_reg[20][2]  ( .D(n3910), .CLK(clk), .Q(\ram[20][2] ) );
  DFFNX1 \ram_reg[20][1]  ( .D(n3909), .CLK(clk), .Q(\ram[20][1] ) );
  DFFNX1 \ram_reg[20][0]  ( .D(n3908), .CLK(clk), .Q(\ram[20][0] ) );
  DFFNX1 \ram_reg[21][7]  ( .D(n3907), .CLK(clk), .Q(\ram[21][7] ) );
  DFFNX1 \ram_reg[21][6]  ( .D(n3906), .CLK(clk), .Q(\ram[21][6] ) );
  DFFNX1 \ram_reg[21][5]  ( .D(n3905), .CLK(clk), .Q(\ram[21][5] ) );
  DFFNX1 \ram_reg[21][4]  ( .D(n3904), .CLK(clk), .Q(\ram[21][4] ) );
  DFFNX1 \ram_reg[21][3]  ( .D(n3903), .CLK(clk), .Q(\ram[21][3] ) );
  DFFNX1 \ram_reg[21][2]  ( .D(n3902), .CLK(clk), .Q(\ram[21][2] ) );
  DFFNX1 \ram_reg[21][1]  ( .D(n3901), .CLK(clk), .Q(\ram[21][1] ) );
  DFFNX1 \ram_reg[21][0]  ( .D(n3900), .CLK(clk), .Q(\ram[21][0] ) );
  DFFNX1 \ram_reg[22][7]  ( .D(n3899), .CLK(clk), .Q(\ram[22][7] ) );
  DFFNX1 \ram_reg[22][6]  ( .D(n3898), .CLK(clk), .Q(\ram[22][6] ) );
  DFFNX1 \ram_reg[22][5]  ( .D(n3897), .CLK(clk), .Q(\ram[22][5] ) );
  DFFNX1 \ram_reg[22][4]  ( .D(n3896), .CLK(clk), .Q(\ram[22][4] ) );
  DFFNX1 \ram_reg[22][3]  ( .D(n3895), .CLK(clk), .Q(\ram[22][3] ) );
  DFFNX1 \ram_reg[22][2]  ( .D(n3894), .CLK(clk), .Q(\ram[22][2] ) );
  DFFNX1 \ram_reg[22][1]  ( .D(n3893), .CLK(clk), .Q(\ram[22][1] ) );
  DFFNX1 \ram_reg[22][0]  ( .D(n3892), .CLK(clk), .Q(\ram[22][0] ) );
  DFFNX1 \ram_reg[23][7]  ( .D(n3891), .CLK(clk), .Q(\ram[23][7] ) );
  DFFNX1 \ram_reg[23][6]  ( .D(n3890), .CLK(clk), .Q(\ram[23][6] ) );
  DFFNX1 \ram_reg[23][5]  ( .D(n3889), .CLK(clk), .Q(\ram[23][5] ) );
  DFFNX1 \ram_reg[23][4]  ( .D(n3888), .CLK(clk), .Q(\ram[23][4] ) );
  DFFNX1 \ram_reg[23][3]  ( .D(n3887), .CLK(clk), .Q(\ram[23][3] ) );
  DFFNX1 \ram_reg[23][2]  ( .D(n3886), .CLK(clk), .Q(\ram[23][2] ) );
  DFFNX1 \ram_reg[23][1]  ( .D(n3885), .CLK(clk), .Q(\ram[23][1] ) );
  DFFNX1 \ram_reg[23][0]  ( .D(n3884), .CLK(clk), .Q(\ram[23][0] ) );
  DFFNX1 \ram_reg[24][7]  ( .D(n3883), .CLK(clk), .Q(\ram[24][7] ) );
  DFFNX1 \ram_reg[24][6]  ( .D(n3882), .CLK(clk), .Q(\ram[24][6] ) );
  DFFNX1 \ram_reg[24][5]  ( .D(n3881), .CLK(clk), .Q(\ram[24][5] ) );
  DFFNX1 \ram_reg[24][4]  ( .D(n3880), .CLK(clk), .Q(\ram[24][4] ) );
  DFFNX1 \ram_reg[24][3]  ( .D(n3879), .CLK(clk), .Q(\ram[24][3] ) );
  DFFNX1 \ram_reg[24][2]  ( .D(n3878), .CLK(clk), .Q(\ram[24][2] ) );
  DFFNX1 \ram_reg[24][1]  ( .D(n3877), .CLK(clk), .Q(\ram[24][1] ) );
  DFFNX1 \ram_reg[24][0]  ( .D(n3876), .CLK(clk), .Q(\ram[24][0] ) );
  DFFNX1 \ram_reg[25][7]  ( .D(n3875), .CLK(clk), .Q(\ram[25][7] ) );
  DFFNX1 \ram_reg[25][6]  ( .D(n3874), .CLK(clk), .Q(\ram[25][6] ) );
  DFFNX1 \ram_reg[25][5]  ( .D(n3873), .CLK(clk), .Q(\ram[25][5] ) );
  DFFNX1 \ram_reg[25][4]  ( .D(n3872), .CLK(clk), .Q(\ram[25][4] ) );
  DFFNX1 \ram_reg[25][3]  ( .D(n3871), .CLK(clk), .Q(\ram[25][3] ) );
  DFFNX1 \ram_reg[25][2]  ( .D(n3870), .CLK(clk), .Q(\ram[25][2] ) );
  DFFNX1 \ram_reg[25][1]  ( .D(n3869), .CLK(clk), .Q(\ram[25][1] ) );
  DFFNX1 \ram_reg[25][0]  ( .D(n3868), .CLK(clk), .Q(\ram[25][0] ) );
  DFFNX1 \ram_reg[26][7]  ( .D(n3867), .CLK(clk), .Q(\ram[26][7] ) );
  DFFNX1 \ram_reg[26][6]  ( .D(n3866), .CLK(clk), .Q(\ram[26][6] ) );
  DFFNX1 \ram_reg[26][5]  ( .D(n3865), .CLK(clk), .Q(\ram[26][5] ) );
  DFFNX1 \ram_reg[26][4]  ( .D(n3864), .CLK(clk), .Q(\ram[26][4] ) );
  DFFNX1 \ram_reg[26][3]  ( .D(n3863), .CLK(clk), .Q(\ram[26][3] ) );
  DFFNX1 \ram_reg[26][2]  ( .D(n3862), .CLK(clk), .Q(\ram[26][2] ) );
  DFFNX1 \ram_reg[26][1]  ( .D(n3861), .CLK(clk), .Q(\ram[26][1] ) );
  DFFNX1 \ram_reg[26][0]  ( .D(n3860), .CLK(clk), .Q(\ram[26][0] ) );
  DFFNX1 \ram_reg[27][7]  ( .D(n3859), .CLK(clk), .Q(\ram[27][7] ) );
  DFFNX1 \ram_reg[27][6]  ( .D(n3858), .CLK(clk), .Q(\ram[27][6] ) );
  DFFNX1 \ram_reg[27][5]  ( .D(n3857), .CLK(clk), .Q(\ram[27][5] ) );
  DFFNX1 \ram_reg[27][4]  ( .D(n3856), .CLK(clk), .Q(\ram[27][4] ) );
  DFFNX1 \ram_reg[27][3]  ( .D(n3855), .CLK(clk), .Q(\ram[27][3] ) );
  DFFNX1 \ram_reg[27][2]  ( .D(n3854), .CLK(clk), .Q(\ram[27][2] ) );
  DFFNX1 \ram_reg[27][1]  ( .D(n3853), .CLK(clk), .Q(\ram[27][1] ) );
  DFFNX1 \ram_reg[27][0]  ( .D(n3852), .CLK(clk), .Q(\ram[27][0] ) );
  DFFNX1 \ram_reg[28][7]  ( .D(n3851), .CLK(clk), .Q(\ram[28][7] ) );
  DFFNX1 \ram_reg[28][6]  ( .D(n3850), .CLK(clk), .Q(\ram[28][6] ) );
  DFFNX1 \ram_reg[28][5]  ( .D(n3849), .CLK(clk), .Q(\ram[28][5] ) );
  DFFNX1 \ram_reg[28][4]  ( .D(n3848), .CLK(clk), .Q(\ram[28][4] ) );
  DFFNX1 \ram_reg[28][3]  ( .D(n3847), .CLK(clk), .Q(\ram[28][3] ) );
  DFFNX1 \ram_reg[28][2]  ( .D(n3846), .CLK(clk), .Q(\ram[28][2] ) );
  DFFNX1 \ram_reg[28][1]  ( .D(n3845), .CLK(clk), .Q(\ram[28][1] ) );
  DFFNX1 \ram_reg[28][0]  ( .D(n3844), .CLK(clk), .Q(\ram[28][0] ) );
  DFFNX1 \ram_reg[29][7]  ( .D(n3843), .CLK(clk), .Q(\ram[29][7] ) );
  DFFNX1 \ram_reg[29][6]  ( .D(n3842), .CLK(clk), .Q(\ram[29][6] ) );
  DFFNX1 \ram_reg[29][5]  ( .D(n3841), .CLK(clk), .Q(\ram[29][5] ) );
  DFFNX1 \ram_reg[29][4]  ( .D(n3840), .CLK(clk), .Q(\ram[29][4] ) );
  DFFNX1 \ram_reg[29][3]  ( .D(n3839), .CLK(clk), .Q(\ram[29][3] ) );
  DFFNX1 \ram_reg[29][2]  ( .D(n3838), .CLK(clk), .Q(\ram[29][2] ) );
  DFFNX1 \ram_reg[29][1]  ( .D(n3837), .CLK(clk), .Q(\ram[29][1] ) );
  DFFNX1 \ram_reg[29][0]  ( .D(n3836), .CLK(clk), .Q(\ram[29][0] ) );
  DFFNX1 \ram_reg[30][7]  ( .D(n3835), .CLK(clk), .Q(\ram[30][7] ) );
  DFFNX1 \ram_reg[30][6]  ( .D(n3834), .CLK(clk), .Q(\ram[30][6] ) );
  DFFNX1 \ram_reg[30][5]  ( .D(n3833), .CLK(clk), .Q(\ram[30][5] ) );
  DFFNX1 \ram_reg[30][4]  ( .D(n3832), .CLK(clk), .Q(\ram[30][4] ) );
  DFFNX1 \ram_reg[30][3]  ( .D(n3831), .CLK(clk), .Q(\ram[30][3] ) );
  DFFNX1 \ram_reg[30][2]  ( .D(n3830), .CLK(clk), .Q(\ram[30][2] ) );
  DFFNX1 \ram_reg[30][1]  ( .D(n3829), .CLK(clk), .Q(\ram[30][1] ) );
  DFFNX1 \ram_reg[30][0]  ( .D(n3828), .CLK(clk), .Q(\ram[30][0] ) );
  DFFNX1 \ram_reg[31][7]  ( .D(n3827), .CLK(clk), .Q(\ram[31][7] ) );
  DFFNX1 \ram_reg[31][6]  ( .D(n3826), .CLK(clk), .Q(\ram[31][6] ) );
  DFFNX1 \ram_reg[31][5]  ( .D(n3825), .CLK(clk), .Q(\ram[31][5] ) );
  DFFNX1 \ram_reg[31][4]  ( .D(n3824), .CLK(clk), .Q(\ram[31][4] ) );
  DFFNX1 \ram_reg[31][3]  ( .D(n3823), .CLK(clk), .Q(\ram[31][3] ) );
  DFFNX1 \ram_reg[31][2]  ( .D(n3822), .CLK(clk), .Q(\ram[31][2] ) );
  DFFNX1 \ram_reg[31][1]  ( .D(n3821), .CLK(clk), .Q(\ram[31][1] ) );
  DFFNX1 \ram_reg[31][0]  ( .D(n3820), .CLK(clk), .Q(\ram[31][0] ) );
  DFFNX1 \ram_reg[32][7]  ( .D(n3819), .CLK(clk), .Q(\ram[32][7] ) );
  DFFNX1 \ram_reg[32][6]  ( .D(n3818), .CLK(clk), .Q(\ram[32][6] ) );
  DFFNX1 \ram_reg[32][5]  ( .D(n3817), .CLK(clk), .Q(\ram[32][5] ) );
  DFFNX1 \ram_reg[32][4]  ( .D(n3816), .CLK(clk), .Q(\ram[32][4] ) );
  DFFNX1 \ram_reg[32][3]  ( .D(n3815), .CLK(clk), .Q(\ram[32][3] ) );
  DFFNX1 \ram_reg[32][2]  ( .D(n3814), .CLK(clk), .Q(\ram[32][2] ) );
  DFFNX1 \ram_reg[32][1]  ( .D(n3813), .CLK(clk), .Q(\ram[32][1] ) );
  DFFNX1 \ram_reg[32][0]  ( .D(n3812), .CLK(clk), .Q(\ram[32][0] ) );
  DFFNX1 \ram_reg[33][7]  ( .D(n3811), .CLK(clk), .Q(\ram[33][7] ) );
  DFFNX1 \ram_reg[33][6]  ( .D(n3810), .CLK(clk), .Q(\ram[33][6] ) );
  DFFNX1 \ram_reg[33][5]  ( .D(n3809), .CLK(clk), .Q(\ram[33][5] ) );
  DFFNX1 \ram_reg[33][4]  ( .D(n3808), .CLK(clk), .Q(\ram[33][4] ) );
  DFFNX1 \ram_reg[33][3]  ( .D(n3807), .CLK(clk), .Q(\ram[33][3] ) );
  DFFNX1 \ram_reg[33][2]  ( .D(n3806), .CLK(clk), .Q(\ram[33][2] ) );
  DFFNX1 \ram_reg[33][1]  ( .D(n3805), .CLK(clk), .Q(\ram[33][1] ) );
  DFFNX1 \ram_reg[33][0]  ( .D(n3804), .CLK(clk), .Q(\ram[33][0] ) );
  DFFNX1 \ram_reg[34][7]  ( .D(n3803), .CLK(clk), .Q(\ram[34][7] ) );
  DFFNX1 \ram_reg[34][6]  ( .D(n3802), .CLK(clk), .Q(\ram[34][6] ) );
  DFFNX1 \ram_reg[34][5]  ( .D(n3801), .CLK(clk), .Q(\ram[34][5] ) );
  DFFNX1 \ram_reg[34][4]  ( .D(n3800), .CLK(clk), .Q(\ram[34][4] ) );
  DFFNX1 \ram_reg[34][3]  ( .D(n3799), .CLK(clk), .Q(\ram[34][3] ) );
  DFFNX1 \ram_reg[34][2]  ( .D(n3798), .CLK(clk), .Q(\ram[34][2] ) );
  DFFNX1 \ram_reg[34][1]  ( .D(n3797), .CLK(clk), .Q(\ram[34][1] ) );
  DFFNX1 \ram_reg[34][0]  ( .D(n3796), .CLK(clk), .Q(\ram[34][0] ) );
  DFFNX1 \ram_reg[35][7]  ( .D(n3795), .CLK(clk), .Q(\ram[35][7] ) );
  DFFNX1 \ram_reg[35][6]  ( .D(n3794), .CLK(clk), .Q(\ram[35][6] ) );
  DFFNX1 \ram_reg[35][5]  ( .D(n3793), .CLK(clk), .Q(\ram[35][5] ) );
  DFFNX1 \ram_reg[35][4]  ( .D(n3792), .CLK(clk), .Q(\ram[35][4] ) );
  DFFNX1 \ram_reg[35][3]  ( .D(n3791), .CLK(clk), .Q(\ram[35][3] ) );
  DFFNX1 \ram_reg[35][2]  ( .D(n3790), .CLK(clk), .Q(\ram[35][2] ) );
  DFFNX1 \ram_reg[35][1]  ( .D(n3789), .CLK(clk), .Q(\ram[35][1] ) );
  DFFNX1 \ram_reg[35][0]  ( .D(n3788), .CLK(clk), .Q(\ram[35][0] ) );
  DFFNX1 \ram_reg[36][7]  ( .D(n3787), .CLK(clk), .Q(\ram[36][7] ) );
  DFFNX1 \ram_reg[36][6]  ( .D(n3786), .CLK(clk), .Q(\ram[36][6] ) );
  DFFNX1 \ram_reg[36][5]  ( .D(n3785), .CLK(clk), .Q(\ram[36][5] ) );
  DFFNX1 \ram_reg[36][4]  ( .D(n3784), .CLK(clk), .Q(\ram[36][4] ) );
  DFFNX1 \ram_reg[36][3]  ( .D(n3783), .CLK(clk), .Q(\ram[36][3] ) );
  DFFNX1 \ram_reg[36][2]  ( .D(n3782), .CLK(clk), .Q(\ram[36][2] ) );
  DFFNX1 \ram_reg[36][1]  ( .D(n3781), .CLK(clk), .Q(\ram[36][1] ) );
  DFFNX1 \ram_reg[36][0]  ( .D(n3780), .CLK(clk), .Q(\ram[36][0] ) );
  DFFNX1 \ram_reg[37][7]  ( .D(n3779), .CLK(clk), .Q(\ram[37][7] ) );
  DFFNX1 \ram_reg[37][6]  ( .D(n3778), .CLK(clk), .Q(\ram[37][6] ) );
  DFFNX1 \ram_reg[37][5]  ( .D(n3777), .CLK(clk), .Q(\ram[37][5] ) );
  DFFNX1 \ram_reg[37][4]  ( .D(n3776), .CLK(clk), .Q(\ram[37][4] ) );
  DFFNX1 \ram_reg[37][3]  ( .D(n3775), .CLK(clk), .Q(\ram[37][3] ) );
  DFFNX1 \ram_reg[37][2]  ( .D(n3774), .CLK(clk), .Q(\ram[37][2] ) );
  DFFNX1 \ram_reg[37][1]  ( .D(n3773), .CLK(clk), .Q(\ram[37][1] ) );
  DFFNX1 \ram_reg[37][0]  ( .D(n3772), .CLK(clk), .Q(\ram[37][0] ) );
  DFFNX1 \ram_reg[38][7]  ( .D(n3771), .CLK(clk), .Q(\ram[38][7] ) );
  DFFNX1 \ram_reg[38][6]  ( .D(n3770), .CLK(clk), .Q(\ram[38][6] ) );
  DFFNX1 \ram_reg[38][5]  ( .D(n3769), .CLK(clk), .Q(\ram[38][5] ) );
  DFFNX1 \ram_reg[38][4]  ( .D(n3768), .CLK(clk), .Q(\ram[38][4] ) );
  DFFNX1 \ram_reg[38][3]  ( .D(n3767), .CLK(clk), .Q(\ram[38][3] ) );
  DFFNX1 \ram_reg[38][2]  ( .D(n3766), .CLK(clk), .Q(\ram[38][2] ) );
  DFFNX1 \ram_reg[38][1]  ( .D(n3765), .CLK(clk), .Q(\ram[38][1] ) );
  DFFNX1 \ram_reg[38][0]  ( .D(n3764), .CLK(clk), .Q(\ram[38][0] ) );
  DFFNX1 \ram_reg[39][7]  ( .D(n3763), .CLK(clk), .Q(\ram[39][7] ) );
  DFFNX1 \ram_reg[39][6]  ( .D(n3762), .CLK(clk), .Q(\ram[39][6] ) );
  DFFNX1 \ram_reg[39][5]  ( .D(n3761), .CLK(clk), .Q(\ram[39][5] ) );
  DFFNX1 \ram_reg[39][4]  ( .D(n3760), .CLK(clk), .Q(\ram[39][4] ) );
  DFFNX1 \ram_reg[39][3]  ( .D(n3759), .CLK(clk), .Q(\ram[39][3] ) );
  DFFNX1 \ram_reg[39][2]  ( .D(n3758), .CLK(clk), .Q(\ram[39][2] ) );
  DFFNX1 \ram_reg[39][1]  ( .D(n3757), .CLK(clk), .Q(\ram[39][1] ) );
  DFFNX1 \ram_reg[39][0]  ( .D(n3756), .CLK(clk), .Q(\ram[39][0] ) );
  DFFNX1 \ram_reg[40][7]  ( .D(n3755), .CLK(clk), .Q(\ram[40][7] ) );
  DFFNX1 \ram_reg[40][6]  ( .D(n3754), .CLK(clk), .Q(\ram[40][6] ) );
  DFFNX1 \ram_reg[40][5]  ( .D(n3753), .CLK(clk), .Q(\ram[40][5] ) );
  DFFNX1 \ram_reg[40][4]  ( .D(n3752), .CLK(clk), .Q(\ram[40][4] ) );
  DFFNX1 \ram_reg[40][3]  ( .D(n3751), .CLK(clk), .Q(\ram[40][3] ) );
  DFFNX1 \ram_reg[40][2]  ( .D(n3750), .CLK(clk), .Q(\ram[40][2] ) );
  DFFNX1 \ram_reg[40][1]  ( .D(n3749), .CLK(clk), .Q(\ram[40][1] ) );
  DFFNX1 \ram_reg[40][0]  ( .D(n3748), .CLK(clk), .Q(\ram[40][0] ) );
  DFFNX1 \ram_reg[41][7]  ( .D(n3747), .CLK(clk), .Q(\ram[41][7] ) );
  DFFNX1 \ram_reg[41][6]  ( .D(n3746), .CLK(clk), .Q(\ram[41][6] ) );
  DFFNX1 \ram_reg[41][5]  ( .D(n3745), .CLK(clk), .Q(\ram[41][5] ) );
  DFFNX1 \ram_reg[41][4]  ( .D(n3744), .CLK(clk), .Q(\ram[41][4] ) );
  DFFNX1 \ram_reg[41][3]  ( .D(n3743), .CLK(clk), .Q(\ram[41][3] ) );
  DFFNX1 \ram_reg[41][2]  ( .D(n3742), .CLK(clk), .Q(\ram[41][2] ) );
  DFFNX1 \ram_reg[41][1]  ( .D(n3741), .CLK(clk), .Q(\ram[41][1] ) );
  DFFNX1 \ram_reg[41][0]  ( .D(n3740), .CLK(clk), .Q(\ram[41][0] ) );
  DFFNX1 \ram_reg[42][7]  ( .D(n3739), .CLK(clk), .Q(\ram[42][7] ) );
  DFFNX1 \ram_reg[42][6]  ( .D(n3738), .CLK(clk), .Q(\ram[42][6] ) );
  DFFNX1 \ram_reg[42][5]  ( .D(n3737), .CLK(clk), .Q(\ram[42][5] ) );
  DFFNX1 \ram_reg[42][4]  ( .D(n3736), .CLK(clk), .Q(\ram[42][4] ) );
  DFFNX1 \ram_reg[42][3]  ( .D(n3735), .CLK(clk), .Q(\ram[42][3] ) );
  DFFNX1 \ram_reg[42][2]  ( .D(n3734), .CLK(clk), .Q(\ram[42][2] ) );
  DFFNX1 \ram_reg[42][1]  ( .D(n3733), .CLK(clk), .Q(\ram[42][1] ) );
  DFFNX1 \ram_reg[42][0]  ( .D(n3732), .CLK(clk), .Q(\ram[42][0] ) );
  DFFNX1 \ram_reg[43][7]  ( .D(n3731), .CLK(clk), .Q(\ram[43][7] ) );
  DFFNX1 \ram_reg[43][6]  ( .D(n3730), .CLK(clk), .Q(\ram[43][6] ) );
  DFFNX1 \ram_reg[43][5]  ( .D(n3729), .CLK(clk), .Q(\ram[43][5] ) );
  DFFNX1 \ram_reg[43][4]  ( .D(n3728), .CLK(clk), .Q(\ram[43][4] ) );
  DFFNX1 \ram_reg[43][3]  ( .D(n3727), .CLK(clk), .Q(\ram[43][3] ) );
  DFFNX1 \ram_reg[43][2]  ( .D(n3726), .CLK(clk), .Q(\ram[43][2] ) );
  DFFNX1 \ram_reg[43][1]  ( .D(n3725), .CLK(clk), .Q(\ram[43][1] ) );
  DFFNX1 \ram_reg[43][0]  ( .D(n3724), .CLK(clk), .Q(\ram[43][0] ) );
  DFFNX1 \ram_reg[44][7]  ( .D(n3723), .CLK(clk), .Q(\ram[44][7] ) );
  DFFNX1 \ram_reg[44][6]  ( .D(n3722), .CLK(clk), .Q(\ram[44][6] ) );
  DFFNX1 \ram_reg[44][5]  ( .D(n3721), .CLK(clk), .Q(\ram[44][5] ) );
  DFFNX1 \ram_reg[44][4]  ( .D(n3720), .CLK(clk), .Q(\ram[44][4] ) );
  DFFNX1 \ram_reg[44][3]  ( .D(n3719), .CLK(clk), .Q(\ram[44][3] ) );
  DFFNX1 \ram_reg[44][2]  ( .D(n3718), .CLK(clk), .Q(\ram[44][2] ) );
  DFFNX1 \ram_reg[44][1]  ( .D(n3717), .CLK(clk), .Q(\ram[44][1] ) );
  DFFNX1 \ram_reg[44][0]  ( .D(n3716), .CLK(clk), .Q(\ram[44][0] ) );
  DFFNX1 \ram_reg[45][7]  ( .D(n3715), .CLK(clk), .Q(\ram[45][7] ) );
  DFFNX1 \ram_reg[45][6]  ( .D(n3714), .CLK(clk), .Q(\ram[45][6] ) );
  DFFNX1 \ram_reg[45][5]  ( .D(n3713), .CLK(clk), .Q(\ram[45][5] ) );
  DFFNX1 \ram_reg[45][4]  ( .D(n3712), .CLK(clk), .Q(\ram[45][4] ) );
  DFFNX1 \ram_reg[45][3]  ( .D(n3711), .CLK(clk), .Q(\ram[45][3] ) );
  DFFNX1 \ram_reg[45][2]  ( .D(n3710), .CLK(clk), .Q(\ram[45][2] ) );
  DFFNX1 \ram_reg[45][1]  ( .D(n3709), .CLK(clk), .Q(\ram[45][1] ) );
  DFFNX1 \ram_reg[45][0]  ( .D(n3708), .CLK(clk), .Q(\ram[45][0] ) );
  DFFNX1 \ram_reg[46][7]  ( .D(n3707), .CLK(clk), .Q(\ram[46][7] ) );
  DFFNX1 \ram_reg[46][6]  ( .D(n3706), .CLK(clk), .Q(\ram[46][6] ) );
  DFFNX1 \ram_reg[46][5]  ( .D(n3705), .CLK(clk), .Q(\ram[46][5] ) );
  DFFNX1 \ram_reg[46][4]  ( .D(n3704), .CLK(clk), .Q(\ram[46][4] ) );
  DFFNX1 \ram_reg[46][3]  ( .D(n3703), .CLK(clk), .Q(\ram[46][3] ) );
  DFFNX1 \ram_reg[46][2]  ( .D(n3702), .CLK(clk), .Q(\ram[46][2] ) );
  DFFNX1 \ram_reg[46][1]  ( .D(n3701), .CLK(clk), .Q(\ram[46][1] ) );
  DFFNX1 \ram_reg[46][0]  ( .D(n3700), .CLK(clk), .Q(\ram[46][0] ) );
  DFFNX1 \ram_reg[47][7]  ( .D(n3699), .CLK(clk), .Q(\ram[47][7] ) );
  DFFNX1 \ram_reg[47][6]  ( .D(n3698), .CLK(clk), .Q(\ram[47][6] ) );
  DFFNX1 \ram_reg[47][5]  ( .D(n3697), .CLK(clk), .Q(\ram[47][5] ) );
  DFFNX1 \ram_reg[47][4]  ( .D(n3696), .CLK(clk), .Q(\ram[47][4] ) );
  DFFNX1 \ram_reg[47][3]  ( .D(n3695), .CLK(clk), .Q(\ram[47][3] ) );
  DFFNX1 \ram_reg[47][2]  ( .D(n3694), .CLK(clk), .Q(\ram[47][2] ) );
  DFFNX1 \ram_reg[47][1]  ( .D(n3693), .CLK(clk), .Q(\ram[47][1] ) );
  DFFNX1 \ram_reg[47][0]  ( .D(n3692), .CLK(clk), .Q(\ram[47][0] ) );
  DFFNX1 \ram_reg[48][7]  ( .D(n3691), .CLK(clk), .Q(\ram[48][7] ) );
  DFFNX1 \ram_reg[48][6]  ( .D(n3690), .CLK(clk), .Q(\ram[48][6] ) );
  DFFNX1 \ram_reg[48][5]  ( .D(n3689), .CLK(clk), .Q(\ram[48][5] ) );
  DFFNX1 \ram_reg[48][4]  ( .D(n3688), .CLK(clk), .Q(\ram[48][4] ) );
  DFFNX1 \ram_reg[48][3]  ( .D(n3687), .CLK(clk), .Q(\ram[48][3] ) );
  DFFNX1 \ram_reg[48][2]  ( .D(n3686), .CLK(clk), .Q(\ram[48][2] ) );
  DFFNX1 \ram_reg[48][1]  ( .D(n3685), .CLK(clk), .Q(\ram[48][1] ) );
  DFFNX1 \ram_reg[48][0]  ( .D(n3684), .CLK(clk), .Q(\ram[48][0] ) );
  DFFNX1 \ram_reg[49][7]  ( .D(n3683), .CLK(clk), .Q(\ram[49][7] ) );
  DFFNX1 \ram_reg[49][6]  ( .D(n3682), .CLK(clk), .Q(\ram[49][6] ) );
  DFFNX1 \ram_reg[49][5]  ( .D(n3681), .CLK(clk), .Q(\ram[49][5] ) );
  DFFNX1 \ram_reg[49][4]  ( .D(n3680), .CLK(clk), .Q(\ram[49][4] ) );
  DFFNX1 \ram_reg[49][3]  ( .D(n3679), .CLK(clk), .Q(\ram[49][3] ) );
  DFFNX1 \ram_reg[49][2]  ( .D(n3678), .CLK(clk), .Q(\ram[49][2] ) );
  DFFNX1 \ram_reg[49][1]  ( .D(n3677), .CLK(clk), .Q(\ram[49][1] ) );
  DFFNX1 \ram_reg[49][0]  ( .D(n3676), .CLK(clk), .Q(\ram[49][0] ) );
  DFFNX1 \ram_reg[50][7]  ( .D(n3675), .CLK(clk), .Q(\ram[50][7] ) );
  DFFNX1 \ram_reg[50][6]  ( .D(n3674), .CLK(clk), .Q(\ram[50][6] ) );
  DFFNX1 \ram_reg[50][5]  ( .D(n3673), .CLK(clk), .Q(\ram[50][5] ) );
  DFFNX1 \ram_reg[50][4]  ( .D(n3672), .CLK(clk), .Q(\ram[50][4] ) );
  DFFNX1 \ram_reg[50][3]  ( .D(n3671), .CLK(clk), .Q(\ram[50][3] ) );
  DFFNX1 \ram_reg[50][2]  ( .D(n3670), .CLK(clk), .Q(\ram[50][2] ) );
  DFFNX1 \ram_reg[50][1]  ( .D(n3669), .CLK(clk), .Q(\ram[50][1] ) );
  DFFNX1 \ram_reg[50][0]  ( .D(n3668), .CLK(clk), .Q(\ram[50][0] ) );
  DFFNX1 \ram_reg[51][7]  ( .D(n3667), .CLK(clk), .Q(\ram[51][7] ) );
  DFFNX1 \ram_reg[51][6]  ( .D(n3666), .CLK(clk), .Q(\ram[51][6] ) );
  DFFNX1 \ram_reg[51][5]  ( .D(n3665), .CLK(clk), .Q(\ram[51][5] ) );
  DFFNX1 \ram_reg[51][4]  ( .D(n3664), .CLK(clk), .Q(\ram[51][4] ) );
  DFFNX1 \ram_reg[51][3]  ( .D(n3663), .CLK(clk), .Q(\ram[51][3] ) );
  DFFNX1 \ram_reg[51][2]  ( .D(n3662), .CLK(clk), .Q(\ram[51][2] ) );
  DFFNX1 \ram_reg[51][1]  ( .D(n3661), .CLK(clk), .Q(\ram[51][1] ) );
  DFFNX1 \ram_reg[51][0]  ( .D(n3660), .CLK(clk), .Q(\ram[51][0] ) );
  DFFNX1 \ram_reg[52][7]  ( .D(n3659), .CLK(clk), .Q(\ram[52][7] ) );
  DFFNX1 \ram_reg[52][6]  ( .D(n3658), .CLK(clk), .Q(\ram[52][6] ) );
  DFFNX1 \ram_reg[52][5]  ( .D(n3657), .CLK(clk), .Q(\ram[52][5] ) );
  DFFNX1 \ram_reg[52][4]  ( .D(n3656), .CLK(clk), .Q(\ram[52][4] ) );
  DFFNX1 \ram_reg[52][3]  ( .D(n3655), .CLK(clk), .Q(\ram[52][3] ) );
  DFFNX1 \ram_reg[52][2]  ( .D(n3654), .CLK(clk), .Q(\ram[52][2] ) );
  DFFNX1 \ram_reg[52][1]  ( .D(n3653), .CLK(clk), .Q(\ram[52][1] ) );
  DFFNX1 \ram_reg[52][0]  ( .D(n3652), .CLK(clk), .Q(\ram[52][0] ) );
  DFFNX1 \ram_reg[53][7]  ( .D(n3651), .CLK(clk), .Q(\ram[53][7] ) );
  DFFNX1 \ram_reg[53][6]  ( .D(n3650), .CLK(clk), .Q(\ram[53][6] ) );
  DFFNX1 \ram_reg[53][5]  ( .D(n3649), .CLK(clk), .Q(\ram[53][5] ) );
  DFFNX1 \ram_reg[53][4]  ( .D(n3648), .CLK(clk), .Q(\ram[53][4] ) );
  DFFNX1 \ram_reg[53][3]  ( .D(n3647), .CLK(clk), .Q(\ram[53][3] ) );
  DFFNX1 \ram_reg[53][2]  ( .D(n3646), .CLK(clk), .Q(\ram[53][2] ) );
  DFFNX1 \ram_reg[53][1]  ( .D(n3645), .CLK(clk), .Q(\ram[53][1] ) );
  DFFNX1 \ram_reg[53][0]  ( .D(n3644), .CLK(clk), .Q(\ram[53][0] ) );
  DFFNX1 \ram_reg[54][7]  ( .D(n3643), .CLK(clk), .Q(\ram[54][7] ) );
  DFFNX1 \ram_reg[54][6]  ( .D(n3642), .CLK(clk), .Q(\ram[54][6] ) );
  DFFNX1 \ram_reg[54][5]  ( .D(n3641), .CLK(clk), .Q(\ram[54][5] ) );
  DFFNX1 \ram_reg[54][4]  ( .D(n3640), .CLK(clk), .Q(\ram[54][4] ) );
  DFFNX1 \ram_reg[54][3]  ( .D(n3639), .CLK(clk), .Q(\ram[54][3] ) );
  DFFNX1 \ram_reg[54][2]  ( .D(n3638), .CLK(clk), .Q(\ram[54][2] ) );
  DFFNX1 \ram_reg[54][1]  ( .D(n3637), .CLK(clk), .Q(\ram[54][1] ) );
  DFFNX1 \ram_reg[54][0]  ( .D(n3636), .CLK(clk), .Q(\ram[54][0] ) );
  DFFNX1 \ram_reg[55][7]  ( .D(n3635), .CLK(clk), .Q(\ram[55][7] ) );
  DFFNX1 \ram_reg[55][6]  ( .D(n3634), .CLK(clk), .Q(\ram[55][6] ) );
  DFFNX1 \ram_reg[55][5]  ( .D(n3633), .CLK(clk), .Q(\ram[55][5] ) );
  DFFNX1 \ram_reg[55][4]  ( .D(n3632), .CLK(clk), .Q(\ram[55][4] ) );
  DFFNX1 \ram_reg[55][3]  ( .D(n3631), .CLK(clk), .Q(\ram[55][3] ) );
  DFFNX1 \ram_reg[55][2]  ( .D(n3630), .CLK(clk), .Q(\ram[55][2] ) );
  DFFNX1 \ram_reg[55][1]  ( .D(n3629), .CLK(clk), .Q(\ram[55][1] ) );
  DFFNX1 \ram_reg[55][0]  ( .D(n3628), .CLK(clk), .Q(\ram[55][0] ) );
  DFFNX1 \ram_reg[56][7]  ( .D(n3627), .CLK(clk), .Q(\ram[56][7] ) );
  DFFNX1 \ram_reg[56][6]  ( .D(n3626), .CLK(clk), .Q(\ram[56][6] ) );
  DFFNX1 \ram_reg[56][5]  ( .D(n3625), .CLK(clk), .Q(\ram[56][5] ) );
  DFFNX1 \ram_reg[56][4]  ( .D(n3624), .CLK(clk), .Q(\ram[56][4] ) );
  DFFNX1 \ram_reg[56][3]  ( .D(n3623), .CLK(clk), .Q(\ram[56][3] ) );
  DFFNX1 \ram_reg[56][2]  ( .D(n3622), .CLK(clk), .Q(\ram[56][2] ) );
  DFFNX1 \ram_reg[56][1]  ( .D(n3621), .CLK(clk), .Q(\ram[56][1] ) );
  DFFNX1 \ram_reg[56][0]  ( .D(n3620), .CLK(clk), .Q(\ram[56][0] ) );
  DFFNX1 \ram_reg[57][7]  ( .D(n3619), .CLK(clk), .Q(\ram[57][7] ) );
  DFFNX1 \ram_reg[57][6]  ( .D(n3618), .CLK(clk), .Q(\ram[57][6] ) );
  DFFNX1 \ram_reg[57][5]  ( .D(n3617), .CLK(clk), .Q(\ram[57][5] ) );
  DFFNX1 \ram_reg[57][4]  ( .D(n3616), .CLK(clk), .Q(\ram[57][4] ) );
  DFFNX1 \ram_reg[57][3]  ( .D(n3615), .CLK(clk), .Q(\ram[57][3] ) );
  DFFNX1 \ram_reg[57][2]  ( .D(n3614), .CLK(clk), .Q(\ram[57][2] ) );
  DFFNX1 \ram_reg[57][1]  ( .D(n3613), .CLK(clk), .Q(\ram[57][1] ) );
  DFFNX1 \ram_reg[57][0]  ( .D(n3612), .CLK(clk), .Q(\ram[57][0] ) );
  DFFNX1 \ram_reg[58][7]  ( .D(n3611), .CLK(clk), .Q(\ram[58][7] ) );
  DFFNX1 \ram_reg[58][6]  ( .D(n3610), .CLK(clk), .Q(\ram[58][6] ) );
  DFFNX1 \ram_reg[58][5]  ( .D(n3609), .CLK(clk), .Q(\ram[58][5] ) );
  DFFNX1 \ram_reg[58][4]  ( .D(n3608), .CLK(clk), .Q(\ram[58][4] ) );
  DFFNX1 \ram_reg[58][3]  ( .D(n3607), .CLK(clk), .Q(\ram[58][3] ) );
  DFFNX1 \ram_reg[58][2]  ( .D(n3606), .CLK(clk), .Q(\ram[58][2] ) );
  DFFNX1 \ram_reg[58][1]  ( .D(n3605), .CLK(clk), .Q(\ram[58][1] ) );
  DFFNX1 \ram_reg[58][0]  ( .D(n3604), .CLK(clk), .Q(\ram[58][0] ) );
  DFFNX1 \ram_reg[59][7]  ( .D(n3603), .CLK(clk), .Q(\ram[59][7] ) );
  DFFNX1 \ram_reg[59][6]  ( .D(n3602), .CLK(clk), .Q(\ram[59][6] ) );
  DFFNX1 \ram_reg[59][5]  ( .D(n3601), .CLK(clk), .Q(\ram[59][5] ) );
  DFFNX1 \ram_reg[59][4]  ( .D(n3600), .CLK(clk), .Q(\ram[59][4] ) );
  DFFNX1 \ram_reg[59][3]  ( .D(n3599), .CLK(clk), .Q(\ram[59][3] ) );
  DFFNX1 \ram_reg[59][2]  ( .D(n3598), .CLK(clk), .Q(\ram[59][2] ) );
  DFFNX1 \ram_reg[59][1]  ( .D(n3597), .CLK(clk), .Q(\ram[59][1] ) );
  DFFNX1 \ram_reg[59][0]  ( .D(n3596), .CLK(clk), .Q(\ram[59][0] ) );
  DFFNX1 \ram_reg[60][7]  ( .D(n3595), .CLK(clk), .Q(\ram[60][7] ) );
  DFFNX1 \ram_reg[60][6]  ( .D(n3594), .CLK(clk), .Q(\ram[60][6] ) );
  DFFNX1 \ram_reg[60][5]  ( .D(n3593), .CLK(clk), .Q(\ram[60][5] ) );
  DFFNX1 \ram_reg[60][4]  ( .D(n3592), .CLK(clk), .Q(\ram[60][4] ) );
  DFFNX1 \ram_reg[60][3]  ( .D(n3591), .CLK(clk), .Q(\ram[60][3] ) );
  DFFNX1 \ram_reg[60][2]  ( .D(n3590), .CLK(clk), .Q(\ram[60][2] ) );
  DFFNX1 \ram_reg[60][1]  ( .D(n3589), .CLK(clk), .Q(\ram[60][1] ) );
  DFFNX1 \ram_reg[60][0]  ( .D(n3588), .CLK(clk), .Q(\ram[60][0] ) );
  DFFNX1 \ram_reg[61][7]  ( .D(n3587), .CLK(clk), .Q(\ram[61][7] ) );
  DFFNX1 \ram_reg[61][6]  ( .D(n3586), .CLK(clk), .Q(\ram[61][6] ) );
  DFFNX1 \ram_reg[61][5]  ( .D(n3585), .CLK(clk), .Q(\ram[61][5] ) );
  DFFNX1 \ram_reg[61][4]  ( .D(n3584), .CLK(clk), .Q(\ram[61][4] ) );
  DFFNX1 \ram_reg[61][3]  ( .D(n3583), .CLK(clk), .Q(\ram[61][3] ) );
  DFFNX1 \ram_reg[61][2]  ( .D(n3582), .CLK(clk), .Q(\ram[61][2] ) );
  DFFNX1 \ram_reg[61][1]  ( .D(n3581), .CLK(clk), .Q(\ram[61][1] ) );
  DFFNX1 \ram_reg[61][0]  ( .D(n3580), .CLK(clk), .Q(\ram[61][0] ) );
  DFFNX1 \ram_reg[62][7]  ( .D(n3579), .CLK(clk), .Q(\ram[62][7] ) );
  DFFNX1 \ram_reg[62][6]  ( .D(n3578), .CLK(clk), .Q(\ram[62][6] ) );
  DFFNX1 \ram_reg[62][5]  ( .D(n3577), .CLK(clk), .Q(\ram[62][5] ) );
  DFFNX1 \ram_reg[62][4]  ( .D(n3576), .CLK(clk), .Q(\ram[62][4] ) );
  DFFNX1 \ram_reg[62][3]  ( .D(n3575), .CLK(clk), .Q(\ram[62][3] ) );
  DFFNX1 \ram_reg[62][2]  ( .D(n3574), .CLK(clk), .Q(\ram[62][2] ) );
  DFFNX1 \ram_reg[62][1]  ( .D(n3573), .CLK(clk), .Q(\ram[62][1] ) );
  DFFNX1 \ram_reg[62][0]  ( .D(n3572), .CLK(clk), .Q(\ram[62][0] ) );
  DFFNX1 \ram_reg[63][7]  ( .D(n3571), .CLK(clk), .Q(\ram[63][7] ) );
  DFFNX1 \ram_reg[63][6]  ( .D(n3570), .CLK(clk), .Q(\ram[63][6] ) );
  DFFNX1 \ram_reg[63][5]  ( .D(n3569), .CLK(clk), .Q(\ram[63][5] ) );
  DFFNX1 \ram_reg[63][4]  ( .D(n3568), .CLK(clk), .Q(\ram[63][4] ) );
  DFFNX1 \ram_reg[63][3]  ( .D(n3567), .CLK(clk), .Q(\ram[63][3] ) );
  DFFNX1 \ram_reg[63][2]  ( .D(n3566), .CLK(clk), .Q(\ram[63][2] ) );
  DFFNX1 \ram_reg[63][1]  ( .D(n3565), .CLK(clk), .Q(\ram[63][1] ) );
  DFFNX1 \ram_reg[63][0]  ( .D(n3564), .CLK(clk), .Q(\ram[63][0] ) );
  DFFNX1 \ram_reg[64][7]  ( .D(n3563), .CLK(clk), .Q(\ram[64][7] ) );
  DFFNX1 \ram_reg[64][6]  ( .D(n3562), .CLK(clk), .Q(\ram[64][6] ) );
  DFFNX1 \ram_reg[64][5]  ( .D(n3561), .CLK(clk), .Q(\ram[64][5] ) );
  DFFNX1 \ram_reg[64][4]  ( .D(n3560), .CLK(clk), .Q(\ram[64][4] ) );
  DFFNX1 \ram_reg[64][3]  ( .D(n3559), .CLK(clk), .Q(\ram[64][3] ) );
  DFFNX1 \ram_reg[64][2]  ( .D(n3558), .CLK(clk), .Q(\ram[64][2] ) );
  DFFNX1 \ram_reg[64][1]  ( .D(n3557), .CLK(clk), .Q(\ram[64][1] ) );
  DFFNX1 \ram_reg[64][0]  ( .D(n3556), .CLK(clk), .Q(\ram[64][0] ) );
  DFFNX1 \ram_reg[65][7]  ( .D(n3555), .CLK(clk), .Q(\ram[65][7] ) );
  DFFNX1 \ram_reg[65][6]  ( .D(n3554), .CLK(clk), .Q(\ram[65][6] ) );
  DFFNX1 \ram_reg[65][5]  ( .D(n3553), .CLK(clk), .Q(\ram[65][5] ) );
  DFFNX1 \ram_reg[65][4]  ( .D(n3552), .CLK(clk), .Q(\ram[65][4] ) );
  DFFNX1 \ram_reg[65][3]  ( .D(n3551), .CLK(clk), .Q(\ram[65][3] ) );
  DFFNX1 \ram_reg[65][2]  ( .D(n3550), .CLK(clk), .Q(\ram[65][2] ) );
  DFFNX1 \ram_reg[65][1]  ( .D(n3549), .CLK(clk), .Q(\ram[65][1] ) );
  DFFNX1 \ram_reg[65][0]  ( .D(n3548), .CLK(clk), .Q(\ram[65][0] ) );
  DFFNX1 \ram_reg[66][7]  ( .D(n3547), .CLK(clk), .Q(\ram[66][7] ) );
  DFFNX1 \ram_reg[66][6]  ( .D(n3546), .CLK(clk), .Q(\ram[66][6] ) );
  DFFNX1 \ram_reg[66][5]  ( .D(n3545), .CLK(clk), .Q(\ram[66][5] ) );
  DFFNX1 \ram_reg[66][4]  ( .D(n3544), .CLK(clk), .Q(\ram[66][4] ) );
  DFFNX1 \ram_reg[66][3]  ( .D(n3543), .CLK(clk), .Q(\ram[66][3] ) );
  DFFNX1 \ram_reg[66][2]  ( .D(n3542), .CLK(clk), .Q(\ram[66][2] ) );
  DFFNX1 \ram_reg[66][1]  ( .D(n3541), .CLK(clk), .Q(\ram[66][1] ) );
  DFFNX1 \ram_reg[66][0]  ( .D(n3540), .CLK(clk), .Q(\ram[66][0] ) );
  DFFNX1 \ram_reg[67][7]  ( .D(n3539), .CLK(clk), .Q(\ram[67][7] ) );
  DFFNX1 \ram_reg[67][6]  ( .D(n3538), .CLK(clk), .Q(\ram[67][6] ) );
  DFFNX1 \ram_reg[67][5]  ( .D(n3537), .CLK(clk), .Q(\ram[67][5] ) );
  DFFNX1 \ram_reg[67][4]  ( .D(n3536), .CLK(clk), .Q(\ram[67][4] ) );
  DFFNX1 \ram_reg[67][3]  ( .D(n3535), .CLK(clk), .Q(\ram[67][3] ) );
  DFFNX1 \ram_reg[67][2]  ( .D(n3534), .CLK(clk), .Q(\ram[67][2] ) );
  DFFNX1 \ram_reg[67][1]  ( .D(n3533), .CLK(clk), .Q(\ram[67][1] ) );
  DFFNX1 \ram_reg[67][0]  ( .D(n3532), .CLK(clk), .Q(\ram[67][0] ) );
  DFFNX1 \ram_reg[68][7]  ( .D(n3531), .CLK(clk), .Q(\ram[68][7] ) );
  DFFNX1 \ram_reg[68][6]  ( .D(n3530), .CLK(clk), .Q(\ram[68][6] ) );
  DFFNX1 \ram_reg[68][5]  ( .D(n3529), .CLK(clk), .Q(\ram[68][5] ) );
  DFFNX1 \ram_reg[68][4]  ( .D(n3528), .CLK(clk), .Q(\ram[68][4] ) );
  DFFNX1 \ram_reg[68][3]  ( .D(n3527), .CLK(clk), .Q(\ram[68][3] ) );
  DFFNX1 \ram_reg[68][2]  ( .D(n3526), .CLK(clk), .Q(\ram[68][2] ) );
  DFFNX1 \ram_reg[68][1]  ( .D(n3525), .CLK(clk), .Q(\ram[68][1] ) );
  DFFNX1 \ram_reg[68][0]  ( .D(n3524), .CLK(clk), .Q(\ram[68][0] ) );
  DFFNX1 \ram_reg[69][7]  ( .D(n3523), .CLK(clk), .Q(\ram[69][7] ) );
  DFFNX1 \ram_reg[69][6]  ( .D(n3522), .CLK(clk), .Q(\ram[69][6] ) );
  DFFNX1 \ram_reg[69][5]  ( .D(n3521), .CLK(clk), .Q(\ram[69][5] ) );
  DFFNX1 \ram_reg[69][4]  ( .D(n3520), .CLK(clk), .Q(\ram[69][4] ) );
  DFFNX1 \ram_reg[69][3]  ( .D(n3519), .CLK(clk), .Q(\ram[69][3] ) );
  DFFNX1 \ram_reg[69][2]  ( .D(n3518), .CLK(clk), .Q(\ram[69][2] ) );
  DFFNX1 \ram_reg[69][1]  ( .D(n3517), .CLK(clk), .Q(\ram[69][1] ) );
  DFFNX1 \ram_reg[69][0]  ( .D(n3516), .CLK(clk), .Q(\ram[69][0] ) );
  DFFNX1 \ram_reg[70][7]  ( .D(n3515), .CLK(clk), .Q(\ram[70][7] ) );
  DFFNX1 \ram_reg[70][6]  ( .D(n3514), .CLK(clk), .Q(\ram[70][6] ) );
  DFFNX1 \ram_reg[70][5]  ( .D(n3513), .CLK(clk), .Q(\ram[70][5] ) );
  DFFNX1 \ram_reg[70][4]  ( .D(n3512), .CLK(clk), .Q(\ram[70][4] ) );
  DFFNX1 \ram_reg[70][3]  ( .D(n3511), .CLK(clk), .Q(\ram[70][3] ) );
  DFFNX1 \ram_reg[70][2]  ( .D(n3510), .CLK(clk), .Q(\ram[70][2] ) );
  DFFNX1 \ram_reg[70][1]  ( .D(n3509), .CLK(clk), .Q(\ram[70][1] ) );
  DFFNX1 \ram_reg[70][0]  ( .D(n3508), .CLK(clk), .Q(\ram[70][0] ) );
  DFFNX1 \ram_reg[71][7]  ( .D(n3507), .CLK(clk), .Q(\ram[71][7] ) );
  DFFNX1 \ram_reg[71][6]  ( .D(n3506), .CLK(clk), .Q(\ram[71][6] ) );
  DFFNX1 \ram_reg[71][5]  ( .D(n3505), .CLK(clk), .Q(\ram[71][5] ) );
  DFFNX1 \ram_reg[71][4]  ( .D(n3504), .CLK(clk), .Q(\ram[71][4] ) );
  DFFNX1 \ram_reg[71][3]  ( .D(n3503), .CLK(clk), .Q(\ram[71][3] ) );
  DFFNX1 \ram_reg[71][2]  ( .D(n3502), .CLK(clk), .Q(\ram[71][2] ) );
  DFFNX1 \ram_reg[71][1]  ( .D(n3501), .CLK(clk), .Q(\ram[71][1] ) );
  DFFNX1 \ram_reg[71][0]  ( .D(n3500), .CLK(clk), .Q(\ram[71][0] ) );
  DFFNX1 \ram_reg[72][7]  ( .D(n3499), .CLK(clk), .Q(\ram[72][7] ) );
  DFFNX1 \ram_reg[72][6]  ( .D(n3498), .CLK(clk), .Q(\ram[72][6] ) );
  DFFNX1 \ram_reg[72][5]  ( .D(n3497), .CLK(clk), .Q(\ram[72][5] ) );
  DFFNX1 \ram_reg[72][4]  ( .D(n3496), .CLK(clk), .Q(\ram[72][4] ) );
  DFFNX1 \ram_reg[72][3]  ( .D(n3495), .CLK(clk), .Q(\ram[72][3] ) );
  DFFNX1 \ram_reg[72][2]  ( .D(n3494), .CLK(clk), .Q(\ram[72][2] ) );
  DFFNX1 \ram_reg[72][1]  ( .D(n3493), .CLK(clk), .Q(\ram[72][1] ) );
  DFFNX1 \ram_reg[72][0]  ( .D(n3492), .CLK(clk), .Q(\ram[72][0] ) );
  DFFNX1 \ram_reg[73][7]  ( .D(n3491), .CLK(clk), .Q(\ram[73][7] ) );
  DFFNX1 \ram_reg[73][6]  ( .D(n3490), .CLK(clk), .Q(\ram[73][6] ) );
  DFFNX1 \ram_reg[73][5]  ( .D(n3489), .CLK(clk), .Q(\ram[73][5] ) );
  DFFNX1 \ram_reg[73][4]  ( .D(n3488), .CLK(clk), .Q(\ram[73][4] ) );
  DFFNX1 \ram_reg[73][3]  ( .D(n3487), .CLK(clk), .Q(\ram[73][3] ) );
  DFFNX1 \ram_reg[73][2]  ( .D(n3486), .CLK(clk), .Q(\ram[73][2] ) );
  DFFNX1 \ram_reg[73][1]  ( .D(n3485), .CLK(clk), .Q(\ram[73][1] ) );
  DFFNX1 \ram_reg[73][0]  ( .D(n3484), .CLK(clk), .Q(\ram[73][0] ) );
  DFFNX1 \ram_reg[74][7]  ( .D(n3483), .CLK(clk), .Q(\ram[74][7] ) );
  DFFNX1 \ram_reg[74][6]  ( .D(n3482), .CLK(clk), .Q(\ram[74][6] ) );
  DFFNX1 \ram_reg[74][5]  ( .D(n3481), .CLK(clk), .Q(\ram[74][5] ) );
  DFFNX1 \ram_reg[74][4]  ( .D(n3480), .CLK(clk), .Q(\ram[74][4] ) );
  DFFNX1 \ram_reg[74][3]  ( .D(n3479), .CLK(clk), .Q(\ram[74][3] ) );
  DFFNX1 \ram_reg[74][2]  ( .D(n3478), .CLK(clk), .Q(\ram[74][2] ) );
  DFFNX1 \ram_reg[74][1]  ( .D(n3477), .CLK(clk), .Q(\ram[74][1] ) );
  DFFNX1 \ram_reg[74][0]  ( .D(n3476), .CLK(clk), .Q(\ram[74][0] ) );
  DFFNX1 \ram_reg[75][7]  ( .D(n3475), .CLK(clk), .Q(\ram[75][7] ) );
  DFFNX1 \ram_reg[75][6]  ( .D(n3474), .CLK(clk), .Q(\ram[75][6] ) );
  DFFNX1 \ram_reg[75][5]  ( .D(n3473), .CLK(clk), .Q(\ram[75][5] ) );
  DFFNX1 \ram_reg[75][4]  ( .D(n3472), .CLK(clk), .Q(\ram[75][4] ) );
  DFFNX1 \ram_reg[75][3]  ( .D(n3471), .CLK(clk), .Q(\ram[75][3] ) );
  DFFNX1 \ram_reg[75][2]  ( .D(n3470), .CLK(clk), .Q(\ram[75][2] ) );
  DFFNX1 \ram_reg[75][1]  ( .D(n3469), .CLK(clk), .Q(\ram[75][1] ) );
  DFFNX1 \ram_reg[75][0]  ( .D(n3468), .CLK(clk), .Q(\ram[75][0] ) );
  DFFNX1 \ram_reg[76][7]  ( .D(n3467), .CLK(clk), .Q(\ram[76][7] ) );
  DFFNX1 \ram_reg[76][6]  ( .D(n3466), .CLK(clk), .Q(\ram[76][6] ) );
  DFFNX1 \ram_reg[76][5]  ( .D(n3465), .CLK(clk), .Q(\ram[76][5] ) );
  DFFNX1 \ram_reg[76][4]  ( .D(n3464), .CLK(clk), .Q(\ram[76][4] ) );
  DFFNX1 \ram_reg[76][3]  ( .D(n3463), .CLK(clk), .Q(\ram[76][3] ) );
  DFFNX1 \ram_reg[76][2]  ( .D(n3462), .CLK(clk), .Q(\ram[76][2] ) );
  DFFNX1 \ram_reg[76][1]  ( .D(n3461), .CLK(clk), .Q(\ram[76][1] ) );
  DFFNX1 \ram_reg[76][0]  ( .D(n3460), .CLK(clk), .Q(\ram[76][0] ) );
  DFFNX1 \ram_reg[77][7]  ( .D(n3459), .CLK(clk), .Q(\ram[77][7] ) );
  DFFNX1 \ram_reg[77][6]  ( .D(n3458), .CLK(clk), .Q(\ram[77][6] ) );
  DFFNX1 \ram_reg[77][5]  ( .D(n3457), .CLK(clk), .Q(\ram[77][5] ) );
  DFFNX1 \ram_reg[77][4]  ( .D(n3456), .CLK(clk), .Q(\ram[77][4] ) );
  DFFNX1 \ram_reg[77][3]  ( .D(n3455), .CLK(clk), .Q(\ram[77][3] ) );
  DFFNX1 \ram_reg[77][2]  ( .D(n3454), .CLK(clk), .Q(\ram[77][2] ) );
  DFFNX1 \ram_reg[77][1]  ( .D(n3453), .CLK(clk), .Q(\ram[77][1] ) );
  DFFNX1 \ram_reg[77][0]  ( .D(n3452), .CLK(clk), .Q(\ram[77][0] ) );
  DFFNX1 \ram_reg[78][7]  ( .D(n3451), .CLK(clk), .Q(\ram[78][7] ) );
  DFFNX1 \ram_reg[78][6]  ( .D(n3450), .CLK(clk), .Q(\ram[78][6] ) );
  DFFNX1 \ram_reg[78][5]  ( .D(n3449), .CLK(clk), .Q(\ram[78][5] ) );
  DFFNX1 \ram_reg[78][4]  ( .D(n3448), .CLK(clk), .Q(\ram[78][4] ) );
  DFFNX1 \ram_reg[78][3]  ( .D(n3447), .CLK(clk), .Q(\ram[78][3] ) );
  DFFNX1 \ram_reg[78][2]  ( .D(n3446), .CLK(clk), .Q(\ram[78][2] ) );
  DFFNX1 \ram_reg[78][1]  ( .D(n3445), .CLK(clk), .Q(\ram[78][1] ) );
  DFFNX1 \ram_reg[78][0]  ( .D(n3444), .CLK(clk), .Q(\ram[78][0] ) );
  DFFNX1 \ram_reg[79][7]  ( .D(n3443), .CLK(clk), .Q(\ram[79][7] ) );
  DFFNX1 \ram_reg[79][6]  ( .D(n3442), .CLK(clk), .Q(\ram[79][6] ) );
  DFFNX1 \ram_reg[79][5]  ( .D(n3441), .CLK(clk), .Q(\ram[79][5] ) );
  DFFNX1 \ram_reg[79][4]  ( .D(n3440), .CLK(clk), .Q(\ram[79][4] ) );
  DFFNX1 \ram_reg[79][3]  ( .D(n3439), .CLK(clk), .Q(\ram[79][3] ) );
  DFFNX1 \ram_reg[79][2]  ( .D(n3438), .CLK(clk), .Q(\ram[79][2] ) );
  DFFNX1 \ram_reg[79][1]  ( .D(n3437), .CLK(clk), .Q(\ram[79][1] ) );
  DFFNX1 \ram_reg[79][0]  ( .D(n3436), .CLK(clk), .Q(\ram[79][0] ) );
  DFFNX1 \ram_reg[80][7]  ( .D(n3435), .CLK(clk), .Q(\ram[80][7] ) );
  DFFNX1 \ram_reg[80][6]  ( .D(n3434), .CLK(clk), .Q(\ram[80][6] ) );
  DFFNX1 \ram_reg[80][5]  ( .D(n3433), .CLK(clk), .Q(\ram[80][5] ) );
  DFFNX1 \ram_reg[80][4]  ( .D(n3432), .CLK(clk), .Q(\ram[80][4] ) );
  DFFNX1 \ram_reg[80][3]  ( .D(n3431), .CLK(clk), .Q(\ram[80][3] ) );
  DFFNX1 \ram_reg[80][2]  ( .D(n3430), .CLK(clk), .Q(\ram[80][2] ) );
  DFFNX1 \ram_reg[80][1]  ( .D(n3429), .CLK(clk), .Q(\ram[80][1] ) );
  DFFNX1 \ram_reg[80][0]  ( .D(n3428), .CLK(clk), .Q(\ram[80][0] ) );
  DFFNX1 \ram_reg[81][7]  ( .D(n3427), .CLK(clk), .Q(\ram[81][7] ) );
  DFFNX1 \ram_reg[81][6]  ( .D(n3426), .CLK(clk), .Q(\ram[81][6] ) );
  DFFNX1 \ram_reg[81][5]  ( .D(n3425), .CLK(clk), .Q(\ram[81][5] ) );
  DFFNX1 \ram_reg[81][4]  ( .D(n3424), .CLK(clk), .Q(\ram[81][4] ) );
  DFFNX1 \ram_reg[81][3]  ( .D(n3423), .CLK(clk), .Q(\ram[81][3] ) );
  DFFNX1 \ram_reg[81][2]  ( .D(n3422), .CLK(clk), .Q(\ram[81][2] ) );
  DFFNX1 \ram_reg[81][1]  ( .D(n3421), .CLK(clk), .Q(\ram[81][1] ) );
  DFFNX1 \ram_reg[81][0]  ( .D(n3420), .CLK(clk), .Q(\ram[81][0] ) );
  DFFNX1 \ram_reg[82][7]  ( .D(n3419), .CLK(clk), .Q(\ram[82][7] ) );
  DFFNX1 \ram_reg[82][6]  ( .D(n3418), .CLK(clk), .Q(\ram[82][6] ) );
  DFFNX1 \ram_reg[82][5]  ( .D(n3417), .CLK(clk), .Q(\ram[82][5] ) );
  DFFNX1 \ram_reg[82][4]  ( .D(n3416), .CLK(clk), .Q(\ram[82][4] ) );
  DFFNX1 \ram_reg[82][3]  ( .D(n3415), .CLK(clk), .Q(\ram[82][3] ) );
  DFFNX1 \ram_reg[82][2]  ( .D(n3414), .CLK(clk), .Q(\ram[82][2] ) );
  DFFNX1 \ram_reg[82][1]  ( .D(n3413), .CLK(clk), .Q(\ram[82][1] ) );
  DFFNX1 \ram_reg[82][0]  ( .D(n3412), .CLK(clk), .Q(\ram[82][0] ) );
  DFFNX1 \ram_reg[83][7]  ( .D(n3411), .CLK(clk), .Q(\ram[83][7] ) );
  DFFNX1 \ram_reg[83][6]  ( .D(n3410), .CLK(clk), .Q(\ram[83][6] ) );
  DFFNX1 \ram_reg[83][5]  ( .D(n3409), .CLK(clk), .Q(\ram[83][5] ) );
  DFFNX1 \ram_reg[83][4]  ( .D(n3408), .CLK(clk), .Q(\ram[83][4] ) );
  DFFNX1 \ram_reg[83][3]  ( .D(n3407), .CLK(clk), .Q(\ram[83][3] ) );
  DFFNX1 \ram_reg[83][2]  ( .D(n3406), .CLK(clk), .Q(\ram[83][2] ) );
  DFFNX1 \ram_reg[83][1]  ( .D(n3405), .CLK(clk), .Q(\ram[83][1] ) );
  DFFNX1 \ram_reg[83][0]  ( .D(n3404), .CLK(clk), .Q(\ram[83][0] ) );
  DFFNX1 \ram_reg[84][7]  ( .D(n3403), .CLK(clk), .Q(\ram[84][7] ) );
  DFFNX1 \ram_reg[84][6]  ( .D(n3402), .CLK(clk), .Q(\ram[84][6] ) );
  DFFNX1 \ram_reg[84][5]  ( .D(n3401), .CLK(clk), .Q(\ram[84][5] ) );
  DFFNX1 \ram_reg[84][4]  ( .D(n3400), .CLK(clk), .Q(\ram[84][4] ) );
  DFFNX1 \ram_reg[84][3]  ( .D(n3399), .CLK(clk), .Q(\ram[84][3] ) );
  DFFNX1 \ram_reg[84][2]  ( .D(n3398), .CLK(clk), .Q(\ram[84][2] ) );
  DFFNX1 \ram_reg[84][1]  ( .D(n3397), .CLK(clk), .Q(\ram[84][1] ) );
  DFFNX1 \ram_reg[84][0]  ( .D(n3396), .CLK(clk), .Q(\ram[84][0] ) );
  DFFNX1 \ram_reg[85][7]  ( .D(n3395), .CLK(clk), .Q(\ram[85][7] ) );
  DFFNX1 \ram_reg[85][6]  ( .D(n3394), .CLK(clk), .Q(\ram[85][6] ) );
  DFFNX1 \ram_reg[85][5]  ( .D(n3393), .CLK(clk), .Q(\ram[85][5] ) );
  DFFNX1 \ram_reg[85][4]  ( .D(n3392), .CLK(clk), .Q(\ram[85][4] ) );
  DFFNX1 \ram_reg[85][3]  ( .D(n3391), .CLK(clk), .Q(\ram[85][3] ) );
  DFFNX1 \ram_reg[85][2]  ( .D(n3390), .CLK(clk), .Q(\ram[85][2] ) );
  DFFNX1 \ram_reg[85][1]  ( .D(n3389), .CLK(clk), .Q(\ram[85][1] ) );
  DFFNX1 \ram_reg[85][0]  ( .D(n3388), .CLK(clk), .Q(\ram[85][0] ) );
  DFFNX1 \ram_reg[86][7]  ( .D(n3387), .CLK(clk), .Q(\ram[86][7] ) );
  DFFNX1 \ram_reg[86][6]  ( .D(n3386), .CLK(clk), .Q(\ram[86][6] ) );
  DFFNX1 \ram_reg[86][5]  ( .D(n3385), .CLK(clk), .Q(\ram[86][5] ) );
  DFFNX1 \ram_reg[86][4]  ( .D(n3384), .CLK(clk), .Q(\ram[86][4] ) );
  DFFNX1 \ram_reg[86][3]  ( .D(n3383), .CLK(clk), .Q(\ram[86][3] ) );
  DFFNX1 \ram_reg[86][2]  ( .D(n3382), .CLK(clk), .Q(\ram[86][2] ) );
  DFFNX1 \ram_reg[86][1]  ( .D(n3381), .CLK(clk), .Q(\ram[86][1] ) );
  DFFNX1 \ram_reg[86][0]  ( .D(n3380), .CLK(clk), .Q(\ram[86][0] ) );
  DFFNX1 \ram_reg[87][7]  ( .D(n3379), .CLK(clk), .Q(\ram[87][7] ) );
  DFFNX1 \ram_reg[87][6]  ( .D(n3378), .CLK(clk), .Q(\ram[87][6] ) );
  DFFNX1 \ram_reg[87][5]  ( .D(n3377), .CLK(clk), .Q(\ram[87][5] ) );
  DFFNX1 \ram_reg[87][4]  ( .D(n3376), .CLK(clk), .Q(\ram[87][4] ) );
  DFFNX1 \ram_reg[87][3]  ( .D(n3375), .CLK(clk), .Q(\ram[87][3] ) );
  DFFNX1 \ram_reg[87][2]  ( .D(n3374), .CLK(clk), .Q(\ram[87][2] ) );
  DFFNX1 \ram_reg[87][1]  ( .D(n3373), .CLK(clk), .Q(\ram[87][1] ) );
  DFFNX1 \ram_reg[87][0]  ( .D(n3372), .CLK(clk), .Q(\ram[87][0] ) );
  DFFNX1 \ram_reg[88][7]  ( .D(n3371), .CLK(clk), .Q(\ram[88][7] ) );
  DFFNX1 \ram_reg[88][6]  ( .D(n3370), .CLK(clk), .Q(\ram[88][6] ) );
  DFFNX1 \ram_reg[88][5]  ( .D(n3369), .CLK(clk), .Q(\ram[88][5] ) );
  DFFNX1 \ram_reg[88][4]  ( .D(n3368), .CLK(clk), .Q(\ram[88][4] ) );
  DFFNX1 \ram_reg[88][3]  ( .D(n3367), .CLK(clk), .Q(\ram[88][3] ) );
  DFFNX1 \ram_reg[88][2]  ( .D(n3366), .CLK(clk), .Q(\ram[88][2] ) );
  DFFNX1 \ram_reg[88][1]  ( .D(n3365), .CLK(clk), .Q(\ram[88][1] ) );
  DFFNX1 \ram_reg[88][0]  ( .D(n3364), .CLK(clk), .Q(\ram[88][0] ) );
  DFFNX1 \ram_reg[89][7]  ( .D(n3363), .CLK(clk), .Q(\ram[89][7] ) );
  DFFNX1 \ram_reg[89][6]  ( .D(n3362), .CLK(clk), .Q(\ram[89][6] ) );
  DFFNX1 \ram_reg[89][5]  ( .D(n3361), .CLK(clk), .Q(\ram[89][5] ) );
  DFFNX1 \ram_reg[89][4]  ( .D(n3360), .CLK(clk), .Q(\ram[89][4] ) );
  DFFNX1 \ram_reg[89][3]  ( .D(n3359), .CLK(clk), .Q(\ram[89][3] ) );
  DFFNX1 \ram_reg[89][2]  ( .D(n3358), .CLK(clk), .Q(\ram[89][2] ) );
  DFFNX1 \ram_reg[89][1]  ( .D(n3357), .CLK(clk), .Q(\ram[89][1] ) );
  DFFNX1 \ram_reg[89][0]  ( .D(n3356), .CLK(clk), .Q(\ram[89][0] ) );
  DFFNX1 \ram_reg[90][7]  ( .D(n3355), .CLK(clk), .Q(\ram[90][7] ) );
  DFFNX1 \ram_reg[90][6]  ( .D(n3354), .CLK(clk), .Q(\ram[90][6] ) );
  DFFNX1 \ram_reg[90][5]  ( .D(n3353), .CLK(clk), .Q(\ram[90][5] ) );
  DFFNX1 \ram_reg[90][4]  ( .D(n3352), .CLK(clk), .Q(\ram[90][4] ) );
  DFFNX1 \ram_reg[90][3]  ( .D(n3351), .CLK(clk), .Q(\ram[90][3] ) );
  DFFNX1 \ram_reg[90][2]  ( .D(n3350), .CLK(clk), .Q(\ram[90][2] ) );
  DFFNX1 \ram_reg[90][1]  ( .D(n3349), .CLK(clk), .Q(\ram[90][1] ) );
  DFFNX1 \ram_reg[90][0]  ( .D(n3348), .CLK(clk), .Q(\ram[90][0] ) );
  DFFNX1 \ram_reg[91][7]  ( .D(n3347), .CLK(clk), .Q(\ram[91][7] ) );
  DFFNX1 \ram_reg[91][6]  ( .D(n3346), .CLK(clk), .Q(\ram[91][6] ) );
  DFFNX1 \ram_reg[91][5]  ( .D(n3345), .CLK(clk), .Q(\ram[91][5] ) );
  DFFNX1 \ram_reg[91][4]  ( .D(n3344), .CLK(clk), .Q(\ram[91][4] ) );
  DFFNX1 \ram_reg[91][3]  ( .D(n3343), .CLK(clk), .Q(\ram[91][3] ) );
  DFFNX1 \ram_reg[91][2]  ( .D(n3342), .CLK(clk), .Q(\ram[91][2] ) );
  DFFNX1 \ram_reg[91][1]  ( .D(n3341), .CLK(clk), .Q(\ram[91][1] ) );
  DFFNX1 \ram_reg[91][0]  ( .D(n3340), .CLK(clk), .Q(\ram[91][0] ) );
  DFFNX1 \ram_reg[92][7]  ( .D(n3339), .CLK(clk), .Q(\ram[92][7] ) );
  DFFNX1 \ram_reg[92][6]  ( .D(n3338), .CLK(clk), .Q(\ram[92][6] ) );
  DFFNX1 \ram_reg[92][5]  ( .D(n3337), .CLK(clk), .Q(\ram[92][5] ) );
  DFFNX1 \ram_reg[92][4]  ( .D(n3336), .CLK(clk), .Q(\ram[92][4] ) );
  DFFNX1 \ram_reg[92][3]  ( .D(n3335), .CLK(clk), .Q(\ram[92][3] ) );
  DFFNX1 \ram_reg[92][2]  ( .D(n3334), .CLK(clk), .Q(\ram[92][2] ) );
  DFFNX1 \ram_reg[92][1]  ( .D(n3333), .CLK(clk), .Q(\ram[92][1] ) );
  DFFNX1 \ram_reg[92][0]  ( .D(n3332), .CLK(clk), .Q(\ram[92][0] ) );
  DFFNX1 \ram_reg[93][7]  ( .D(n3331), .CLK(clk), .Q(\ram[93][7] ) );
  DFFNX1 \ram_reg[93][6]  ( .D(n3330), .CLK(clk), .Q(\ram[93][6] ) );
  DFFNX1 \ram_reg[93][5]  ( .D(n3329), .CLK(clk), .Q(\ram[93][5] ) );
  DFFNX1 \ram_reg[93][4]  ( .D(n3328), .CLK(clk), .Q(\ram[93][4] ) );
  DFFNX1 \ram_reg[93][3]  ( .D(n3327), .CLK(clk), .Q(\ram[93][3] ) );
  DFFNX1 \ram_reg[93][2]  ( .D(n3326), .CLK(clk), .Q(\ram[93][2] ) );
  DFFNX1 \ram_reg[93][1]  ( .D(n3325), .CLK(clk), .Q(\ram[93][1] ) );
  DFFNX1 \ram_reg[93][0]  ( .D(n3324), .CLK(clk), .Q(\ram[93][0] ) );
  DFFNX1 \ram_reg[94][7]  ( .D(n3323), .CLK(clk), .Q(\ram[94][7] ) );
  DFFNX1 \ram_reg[94][6]  ( .D(n3322), .CLK(clk), .Q(\ram[94][6] ) );
  DFFNX1 \ram_reg[94][5]  ( .D(n3321), .CLK(clk), .Q(\ram[94][5] ) );
  DFFNX1 \ram_reg[94][4]  ( .D(n3320), .CLK(clk), .Q(\ram[94][4] ) );
  DFFNX1 \ram_reg[94][3]  ( .D(n3319), .CLK(clk), .Q(\ram[94][3] ) );
  DFFNX1 \ram_reg[94][2]  ( .D(n3318), .CLK(clk), .Q(\ram[94][2] ) );
  DFFNX1 \ram_reg[94][1]  ( .D(n3317), .CLK(clk), .Q(\ram[94][1] ) );
  DFFNX1 \ram_reg[94][0]  ( .D(n3316), .CLK(clk), .Q(\ram[94][0] ) );
  DFFNX1 \ram_reg[95][7]  ( .D(n3315), .CLK(clk), .Q(\ram[95][7] ) );
  DFFNX1 \ram_reg[95][6]  ( .D(n3314), .CLK(clk), .Q(\ram[95][6] ) );
  DFFNX1 \ram_reg[95][5]  ( .D(n3313), .CLK(clk), .Q(\ram[95][5] ) );
  DFFNX1 \ram_reg[95][4]  ( .D(n3312), .CLK(clk), .Q(\ram[95][4] ) );
  DFFNX1 \ram_reg[95][3]  ( .D(n3311), .CLK(clk), .Q(\ram[95][3] ) );
  DFFNX1 \ram_reg[95][2]  ( .D(n3310), .CLK(clk), .Q(\ram[95][2] ) );
  DFFNX1 \ram_reg[95][1]  ( .D(n3309), .CLK(clk), .Q(\ram[95][1] ) );
  DFFNX1 \ram_reg[95][0]  ( .D(n3308), .CLK(clk), .Q(\ram[95][0] ) );
  DFFNX1 \ram_reg[96][7]  ( .D(n3307), .CLK(clk), .Q(\ram[96][7] ) );
  DFFNX1 \ram_reg[96][6]  ( .D(n3306), .CLK(clk), .Q(\ram[96][6] ) );
  DFFNX1 \ram_reg[96][5]  ( .D(n3305), .CLK(clk), .Q(\ram[96][5] ) );
  DFFNX1 \ram_reg[96][4]  ( .D(n3304), .CLK(clk), .Q(\ram[96][4] ) );
  DFFNX1 \ram_reg[96][3]  ( .D(n3303), .CLK(clk), .Q(\ram[96][3] ) );
  DFFNX1 \ram_reg[96][2]  ( .D(n3302), .CLK(clk), .Q(\ram[96][2] ) );
  DFFNX1 \ram_reg[96][1]  ( .D(n3301), .CLK(clk), .Q(\ram[96][1] ) );
  DFFNX1 \ram_reg[96][0]  ( .D(n3300), .CLK(clk), .Q(\ram[96][0] ) );
  DFFNX1 \ram_reg[97][7]  ( .D(n3299), .CLK(clk), .Q(\ram[97][7] ) );
  DFFNX1 \ram_reg[97][6]  ( .D(n3298), .CLK(clk), .Q(\ram[97][6] ) );
  DFFNX1 \ram_reg[97][5]  ( .D(n3297), .CLK(clk), .Q(\ram[97][5] ) );
  DFFNX1 \ram_reg[97][4]  ( .D(n3296), .CLK(clk), .Q(\ram[97][4] ) );
  DFFNX1 \ram_reg[97][3]  ( .D(n3295), .CLK(clk), .Q(\ram[97][3] ) );
  DFFNX1 \ram_reg[97][2]  ( .D(n3294), .CLK(clk), .Q(\ram[97][2] ) );
  DFFNX1 \ram_reg[97][1]  ( .D(n3293), .CLK(clk), .Q(\ram[97][1] ) );
  DFFNX1 \ram_reg[97][0]  ( .D(n3292), .CLK(clk), .Q(\ram[97][0] ) );
  DFFNX1 \ram_reg[98][7]  ( .D(n3291), .CLK(clk), .Q(\ram[98][7] ) );
  DFFNX1 \ram_reg[98][6]  ( .D(n3290), .CLK(clk), .Q(\ram[98][6] ) );
  DFFNX1 \ram_reg[98][5]  ( .D(n3289), .CLK(clk), .Q(\ram[98][5] ) );
  DFFNX1 \ram_reg[98][4]  ( .D(n3288), .CLK(clk), .Q(\ram[98][4] ) );
  DFFNX1 \ram_reg[98][3]  ( .D(n3287), .CLK(clk), .Q(\ram[98][3] ) );
  DFFNX1 \ram_reg[98][2]  ( .D(n3286), .CLK(clk), .Q(\ram[98][2] ) );
  DFFNX1 \ram_reg[98][1]  ( .D(n3285), .CLK(clk), .Q(\ram[98][1] ) );
  DFFNX1 \ram_reg[98][0]  ( .D(n3284), .CLK(clk), .Q(\ram[98][0] ) );
  DFFNX1 \ram_reg[99][7]  ( .D(n3283), .CLK(clk), .Q(\ram[99][7] ) );
  DFFNX1 \ram_reg[99][6]  ( .D(n3282), .CLK(clk), .Q(\ram[99][6] ) );
  DFFNX1 \ram_reg[99][5]  ( .D(n3281), .CLK(clk), .Q(\ram[99][5] ) );
  DFFNX1 \ram_reg[99][4]  ( .D(n3280), .CLK(clk), .Q(\ram[99][4] ) );
  DFFNX1 \ram_reg[99][3]  ( .D(n3279), .CLK(clk), .Q(\ram[99][3] ) );
  DFFNX1 \ram_reg[99][2]  ( .D(n3278), .CLK(clk), .Q(\ram[99][2] ) );
  DFFNX1 \ram_reg[99][1]  ( .D(n3277), .CLK(clk), .Q(\ram[99][1] ) );
  DFFNX1 \ram_reg[99][0]  ( .D(n3276), .CLK(clk), .Q(\ram[99][0] ) );
  DFFNX1 \ram_reg[100][7]  ( .D(n3275), .CLK(clk), .Q(\ram[100][7] ) );
  DFFNX1 \ram_reg[100][6]  ( .D(n3274), .CLK(clk), .Q(\ram[100][6] ) );
  DFFNX1 \ram_reg[100][5]  ( .D(n3273), .CLK(clk), .Q(\ram[100][5] ) );
  DFFNX1 \ram_reg[100][4]  ( .D(n3272), .CLK(clk), .Q(\ram[100][4] ) );
  DFFNX1 \ram_reg[100][3]  ( .D(n3271), .CLK(clk), .Q(\ram[100][3] ) );
  DFFNX1 \ram_reg[100][2]  ( .D(n3270), .CLK(clk), .Q(\ram[100][2] ) );
  DFFNX1 \ram_reg[100][1]  ( .D(n3269), .CLK(clk), .Q(\ram[100][1] ) );
  DFFNX1 \ram_reg[100][0]  ( .D(n3268), .CLK(clk), .Q(\ram[100][0] ) );
  DFFNX1 \ram_reg[101][7]  ( .D(n3267), .CLK(clk), .Q(\ram[101][7] ) );
  DFFNX1 \ram_reg[101][6]  ( .D(n3266), .CLK(clk), .Q(\ram[101][6] ) );
  DFFNX1 \ram_reg[101][5]  ( .D(n3265), .CLK(clk), .Q(\ram[101][5] ) );
  DFFNX1 \ram_reg[101][4]  ( .D(n3264), .CLK(clk), .Q(\ram[101][4] ) );
  DFFNX1 \ram_reg[101][3]  ( .D(n3263), .CLK(clk), .Q(\ram[101][3] ) );
  DFFNX1 \ram_reg[101][2]  ( .D(n3262), .CLK(clk), .Q(\ram[101][2] ) );
  DFFNX1 \ram_reg[101][1]  ( .D(n3261), .CLK(clk), .Q(\ram[101][1] ) );
  DFFNX1 \ram_reg[101][0]  ( .D(n3260), .CLK(clk), .Q(\ram[101][0] ) );
  DFFNX1 \ram_reg[102][7]  ( .D(n3259), .CLK(clk), .Q(\ram[102][7] ) );
  DFFNX1 \ram_reg[102][6]  ( .D(n3258), .CLK(clk), .Q(\ram[102][6] ) );
  DFFNX1 \ram_reg[102][5]  ( .D(n3257), .CLK(clk), .Q(\ram[102][5] ) );
  DFFNX1 \ram_reg[102][4]  ( .D(n3256), .CLK(clk), .Q(\ram[102][4] ) );
  DFFNX1 \ram_reg[102][3]  ( .D(n3255), .CLK(clk), .Q(\ram[102][3] ) );
  DFFNX1 \ram_reg[102][2]  ( .D(n3254), .CLK(clk), .Q(\ram[102][2] ) );
  DFFNX1 \ram_reg[102][1]  ( .D(n3253), .CLK(clk), .Q(\ram[102][1] ) );
  DFFNX1 \ram_reg[102][0]  ( .D(n3252), .CLK(clk), .Q(\ram[102][0] ) );
  DFFNX1 \ram_reg[103][7]  ( .D(n3251), .CLK(clk), .Q(\ram[103][7] ) );
  DFFNX1 \ram_reg[103][6]  ( .D(n3250), .CLK(clk), .Q(\ram[103][6] ) );
  DFFNX1 \ram_reg[103][5]  ( .D(n3249), .CLK(clk), .Q(\ram[103][5] ) );
  DFFNX1 \ram_reg[103][4]  ( .D(n3248), .CLK(clk), .Q(\ram[103][4] ) );
  DFFNX1 \ram_reg[103][3]  ( .D(n3247), .CLK(clk), .Q(\ram[103][3] ) );
  DFFNX1 \ram_reg[103][2]  ( .D(n3246), .CLK(clk), .Q(\ram[103][2] ) );
  DFFNX1 \ram_reg[103][1]  ( .D(n3245), .CLK(clk), .Q(\ram[103][1] ) );
  DFFNX1 \ram_reg[103][0]  ( .D(n3244), .CLK(clk), .Q(\ram[103][0] ) );
  DFFNX1 \ram_reg[104][7]  ( .D(n3243), .CLK(clk), .Q(\ram[104][7] ) );
  DFFNX1 \ram_reg[104][6]  ( .D(n3242), .CLK(clk), .Q(\ram[104][6] ) );
  DFFNX1 \ram_reg[104][5]  ( .D(n3241), .CLK(clk), .Q(\ram[104][5] ) );
  DFFNX1 \ram_reg[104][4]  ( .D(n3240), .CLK(clk), .Q(\ram[104][4] ) );
  DFFNX1 \ram_reg[104][3]  ( .D(n3239), .CLK(clk), .Q(\ram[104][3] ) );
  DFFNX1 \ram_reg[104][2]  ( .D(n3238), .CLK(clk), .Q(\ram[104][2] ) );
  DFFNX1 \ram_reg[104][1]  ( .D(n3237), .CLK(clk), .Q(\ram[104][1] ) );
  DFFNX1 \ram_reg[104][0]  ( .D(n3236), .CLK(clk), .Q(\ram[104][0] ) );
  DFFNX1 \ram_reg[105][7]  ( .D(n3235), .CLK(clk), .Q(\ram[105][7] ) );
  DFFNX1 \ram_reg[105][6]  ( .D(n3234), .CLK(clk), .Q(\ram[105][6] ) );
  DFFNX1 \ram_reg[105][5]  ( .D(n3233), .CLK(clk), .Q(\ram[105][5] ) );
  DFFNX1 \ram_reg[105][4]  ( .D(n3232), .CLK(clk), .Q(\ram[105][4] ) );
  DFFNX1 \ram_reg[105][3]  ( .D(n3231), .CLK(clk), .Q(\ram[105][3] ) );
  DFFNX1 \ram_reg[105][2]  ( .D(n3230), .CLK(clk), .Q(\ram[105][2] ) );
  DFFNX1 \ram_reg[105][1]  ( .D(n3229), .CLK(clk), .Q(\ram[105][1] ) );
  DFFNX1 \ram_reg[105][0]  ( .D(n3228), .CLK(clk), .Q(\ram[105][0] ) );
  DFFNX1 \ram_reg[106][7]  ( .D(n3227), .CLK(clk), .Q(\ram[106][7] ) );
  DFFNX1 \ram_reg[106][6]  ( .D(n3226), .CLK(clk), .Q(\ram[106][6] ) );
  DFFNX1 \ram_reg[106][5]  ( .D(n3225), .CLK(clk), .Q(\ram[106][5] ) );
  DFFNX1 \ram_reg[106][4]  ( .D(n3224), .CLK(clk), .Q(\ram[106][4] ) );
  DFFNX1 \ram_reg[106][3]  ( .D(n3223), .CLK(clk), .Q(\ram[106][3] ) );
  DFFNX1 \ram_reg[106][2]  ( .D(n3222), .CLK(clk), .Q(\ram[106][2] ) );
  DFFNX1 \ram_reg[106][1]  ( .D(n3221), .CLK(clk), .Q(\ram[106][1] ) );
  DFFNX1 \ram_reg[106][0]  ( .D(n3220), .CLK(clk), .Q(\ram[106][0] ) );
  DFFNX1 \ram_reg[107][7]  ( .D(n3219), .CLK(clk), .Q(\ram[107][7] ) );
  DFFNX1 \ram_reg[107][6]  ( .D(n3218), .CLK(clk), .Q(\ram[107][6] ) );
  DFFNX1 \ram_reg[107][5]  ( .D(n3217), .CLK(clk), .Q(\ram[107][5] ) );
  DFFNX1 \ram_reg[107][4]  ( .D(n3216), .CLK(clk), .Q(\ram[107][4] ) );
  DFFNX1 \ram_reg[107][3]  ( .D(n3215), .CLK(clk), .Q(\ram[107][3] ) );
  DFFNX1 \ram_reg[107][2]  ( .D(n3214), .CLK(clk), .Q(\ram[107][2] ) );
  DFFNX1 \ram_reg[107][1]  ( .D(n3213), .CLK(clk), .Q(\ram[107][1] ) );
  DFFNX1 \ram_reg[107][0]  ( .D(n3212), .CLK(clk), .Q(\ram[107][0] ) );
  DFFNX1 \ram_reg[108][7]  ( .D(n3211), .CLK(clk), .Q(\ram[108][7] ) );
  DFFNX1 \ram_reg[108][6]  ( .D(n3210), .CLK(clk), .Q(\ram[108][6] ) );
  DFFNX1 \ram_reg[108][5]  ( .D(n3209), .CLK(clk), .Q(\ram[108][5] ) );
  DFFNX1 \ram_reg[108][4]  ( .D(n3208), .CLK(clk), .Q(\ram[108][4] ) );
  DFFNX1 \ram_reg[108][3]  ( .D(n3207), .CLK(clk), .Q(\ram[108][3] ) );
  DFFNX1 \ram_reg[108][2]  ( .D(n3206), .CLK(clk), .Q(\ram[108][2] ) );
  DFFNX1 \ram_reg[108][1]  ( .D(n3205), .CLK(clk), .Q(\ram[108][1] ) );
  DFFNX1 \ram_reg[108][0]  ( .D(n3204), .CLK(clk), .Q(\ram[108][0] ) );
  DFFNX1 \ram_reg[109][7]  ( .D(n3203), .CLK(clk), .Q(\ram[109][7] ) );
  DFFNX1 \ram_reg[109][6]  ( .D(n3202), .CLK(clk), .Q(\ram[109][6] ) );
  DFFNX1 \ram_reg[109][5]  ( .D(n3201), .CLK(clk), .Q(\ram[109][5] ) );
  DFFNX1 \ram_reg[109][4]  ( .D(n3200), .CLK(clk), .Q(\ram[109][4] ) );
  DFFNX1 \ram_reg[109][3]  ( .D(n3199), .CLK(clk), .Q(\ram[109][3] ) );
  DFFNX1 \ram_reg[109][2]  ( .D(n3198), .CLK(clk), .Q(\ram[109][2] ) );
  DFFNX1 \ram_reg[109][1]  ( .D(n3197), .CLK(clk), .Q(\ram[109][1] ) );
  DFFNX1 \ram_reg[109][0]  ( .D(n3196), .CLK(clk), .Q(\ram[109][0] ) );
  DFFNX1 \ram_reg[110][7]  ( .D(n3195), .CLK(clk), .Q(\ram[110][7] ) );
  DFFNX1 \ram_reg[110][6]  ( .D(n3194), .CLK(clk), .Q(\ram[110][6] ) );
  DFFNX1 \ram_reg[110][5]  ( .D(n3193), .CLK(clk), .Q(\ram[110][5] ) );
  DFFNX1 \ram_reg[110][4]  ( .D(n3192), .CLK(clk), .Q(\ram[110][4] ) );
  DFFNX1 \ram_reg[110][3]  ( .D(n3191), .CLK(clk), .Q(\ram[110][3] ) );
  DFFNX1 \ram_reg[110][2]  ( .D(n3190), .CLK(clk), .Q(\ram[110][2] ) );
  DFFNX1 \ram_reg[110][1]  ( .D(n3189), .CLK(clk), .Q(\ram[110][1] ) );
  DFFNX1 \ram_reg[110][0]  ( .D(n3188), .CLK(clk), .Q(\ram[110][0] ) );
  DFFNX1 \ram_reg[111][7]  ( .D(n3187), .CLK(clk), .Q(\ram[111][7] ) );
  DFFNX1 \ram_reg[111][6]  ( .D(n3186), .CLK(clk), .Q(\ram[111][6] ) );
  DFFNX1 \ram_reg[111][5]  ( .D(n3185), .CLK(clk), .Q(\ram[111][5] ) );
  DFFNX1 \ram_reg[111][4]  ( .D(n3184), .CLK(clk), .Q(\ram[111][4] ) );
  DFFNX1 \ram_reg[111][3]  ( .D(n3183), .CLK(clk), .Q(\ram[111][3] ) );
  DFFNX1 \ram_reg[111][2]  ( .D(n3182), .CLK(clk), .Q(\ram[111][2] ) );
  DFFNX1 \ram_reg[111][1]  ( .D(n3181), .CLK(clk), .Q(\ram[111][1] ) );
  DFFNX1 \ram_reg[111][0]  ( .D(n3180), .CLK(clk), .Q(\ram[111][0] ) );
  DFFNX1 \ram_reg[112][7]  ( .D(n3179), .CLK(clk), .Q(\ram[112][7] ) );
  DFFNX1 \ram_reg[112][6]  ( .D(n3178), .CLK(clk), .Q(\ram[112][6] ) );
  DFFNX1 \ram_reg[112][5]  ( .D(n3177), .CLK(clk), .Q(\ram[112][5] ) );
  DFFNX1 \ram_reg[112][4]  ( .D(n3176), .CLK(clk), .Q(\ram[112][4] ) );
  DFFNX1 \ram_reg[112][3]  ( .D(n3175), .CLK(clk), .Q(\ram[112][3] ) );
  DFFNX1 \ram_reg[112][2]  ( .D(n3174), .CLK(clk), .Q(\ram[112][2] ) );
  DFFNX1 \ram_reg[112][1]  ( .D(n3173), .CLK(clk), .Q(\ram[112][1] ) );
  DFFNX1 \ram_reg[112][0]  ( .D(n3172), .CLK(clk), .Q(\ram[112][0] ) );
  DFFNX1 \ram_reg[113][7]  ( .D(n3171), .CLK(clk), .Q(\ram[113][7] ) );
  DFFNX1 \ram_reg[113][6]  ( .D(n3170), .CLK(clk), .Q(\ram[113][6] ) );
  DFFNX1 \ram_reg[113][5]  ( .D(n3169), .CLK(clk), .Q(\ram[113][5] ) );
  DFFNX1 \ram_reg[113][4]  ( .D(n3168), .CLK(clk), .Q(\ram[113][4] ) );
  DFFNX1 \ram_reg[113][3]  ( .D(n3167), .CLK(clk), .Q(\ram[113][3] ) );
  DFFNX1 \ram_reg[113][2]  ( .D(n3166), .CLK(clk), .Q(\ram[113][2] ) );
  DFFNX1 \ram_reg[113][1]  ( .D(n3165), .CLK(clk), .Q(\ram[113][1] ) );
  DFFNX1 \ram_reg[113][0]  ( .D(n3164), .CLK(clk), .Q(\ram[113][0] ) );
  DFFNX1 \ram_reg[114][7]  ( .D(n3163), .CLK(clk), .Q(\ram[114][7] ) );
  DFFNX1 \ram_reg[114][6]  ( .D(n3162), .CLK(clk), .Q(\ram[114][6] ) );
  DFFNX1 \ram_reg[114][5]  ( .D(n3161), .CLK(clk), .Q(\ram[114][5] ) );
  DFFNX1 \ram_reg[114][4]  ( .D(n3160), .CLK(clk), .Q(\ram[114][4] ) );
  DFFNX1 \ram_reg[114][3]  ( .D(n3159), .CLK(clk), .Q(\ram[114][3] ) );
  DFFNX1 \ram_reg[114][2]  ( .D(n3158), .CLK(clk), .Q(\ram[114][2] ) );
  DFFNX1 \ram_reg[114][1]  ( .D(n3157), .CLK(clk), .Q(\ram[114][1] ) );
  DFFNX1 \ram_reg[114][0]  ( .D(n3156), .CLK(clk), .Q(\ram[114][0] ) );
  DFFNX1 \ram_reg[115][7]  ( .D(n3155), .CLK(clk), .Q(\ram[115][7] ) );
  DFFNX1 \ram_reg[115][6]  ( .D(n3154), .CLK(clk), .Q(\ram[115][6] ) );
  DFFNX1 \ram_reg[115][5]  ( .D(n3153), .CLK(clk), .Q(\ram[115][5] ) );
  DFFNX1 \ram_reg[115][4]  ( .D(n3152), .CLK(clk), .Q(\ram[115][4] ) );
  DFFNX1 \ram_reg[115][3]  ( .D(n3151), .CLK(clk), .Q(\ram[115][3] ) );
  DFFNX1 \ram_reg[115][2]  ( .D(n3150), .CLK(clk), .Q(\ram[115][2] ) );
  DFFNX1 \ram_reg[115][1]  ( .D(n3149), .CLK(clk), .Q(\ram[115][1] ) );
  DFFNX1 \ram_reg[115][0]  ( .D(n3148), .CLK(clk), .Q(\ram[115][0] ) );
  DFFNX1 \ram_reg[116][7]  ( .D(n3147), .CLK(clk), .Q(\ram[116][7] ) );
  DFFNX1 \ram_reg[116][6]  ( .D(n3146), .CLK(clk), .Q(\ram[116][6] ) );
  DFFNX1 \ram_reg[116][5]  ( .D(n3145), .CLK(clk), .Q(\ram[116][5] ) );
  DFFNX1 \ram_reg[116][4]  ( .D(n3144), .CLK(clk), .Q(\ram[116][4] ) );
  DFFNX1 \ram_reg[116][3]  ( .D(n3143), .CLK(clk), .Q(\ram[116][3] ) );
  DFFNX1 \ram_reg[116][2]  ( .D(n3142), .CLK(clk), .Q(\ram[116][2] ) );
  DFFNX1 \ram_reg[116][1]  ( .D(n3141), .CLK(clk), .Q(\ram[116][1] ) );
  DFFNX1 \ram_reg[116][0]  ( .D(n3140), .CLK(clk), .Q(\ram[116][0] ) );
  DFFNX1 \ram_reg[117][7]  ( .D(n3139), .CLK(clk), .Q(\ram[117][7] ) );
  DFFNX1 \ram_reg[117][6]  ( .D(n3138), .CLK(clk), .Q(\ram[117][6] ) );
  DFFNX1 \ram_reg[117][5]  ( .D(n3137), .CLK(clk), .Q(\ram[117][5] ) );
  DFFNX1 \ram_reg[117][4]  ( .D(n3136), .CLK(clk), .Q(\ram[117][4] ) );
  DFFNX1 \ram_reg[117][3]  ( .D(n3135), .CLK(clk), .Q(\ram[117][3] ) );
  DFFNX1 \ram_reg[117][2]  ( .D(n3134), .CLK(clk), .Q(\ram[117][2] ) );
  DFFNX1 \ram_reg[117][1]  ( .D(n3133), .CLK(clk), .Q(\ram[117][1] ) );
  DFFNX1 \ram_reg[117][0]  ( .D(n3132), .CLK(clk), .Q(\ram[117][0] ) );
  DFFNX1 \ram_reg[118][7]  ( .D(n3131), .CLK(clk), .Q(\ram[118][7] ) );
  DFFNX1 \ram_reg[118][6]  ( .D(n3130), .CLK(clk), .Q(\ram[118][6] ) );
  DFFNX1 \ram_reg[118][5]  ( .D(n3129), .CLK(clk), .Q(\ram[118][5] ) );
  DFFNX1 \ram_reg[118][4]  ( .D(n3128), .CLK(clk), .Q(\ram[118][4] ) );
  DFFNX1 \ram_reg[118][3]  ( .D(n3127), .CLK(clk), .Q(\ram[118][3] ) );
  DFFNX1 \ram_reg[118][2]  ( .D(n3126), .CLK(clk), .Q(\ram[118][2] ) );
  DFFNX1 \ram_reg[118][1]  ( .D(n3125), .CLK(clk), .Q(\ram[118][1] ) );
  DFFNX1 \ram_reg[118][0]  ( .D(n3124), .CLK(clk), .Q(\ram[118][0] ) );
  DFFNX1 \ram_reg[119][7]  ( .D(n3123), .CLK(clk), .Q(\ram[119][7] ) );
  DFFNX1 \ram_reg[119][6]  ( .D(n3122), .CLK(clk), .Q(\ram[119][6] ) );
  DFFNX1 \ram_reg[119][5]  ( .D(n3121), .CLK(clk), .Q(\ram[119][5] ) );
  DFFNX1 \ram_reg[119][4]  ( .D(n3120), .CLK(clk), .Q(\ram[119][4] ) );
  DFFNX1 \ram_reg[119][3]  ( .D(n3119), .CLK(clk), .Q(\ram[119][3] ) );
  DFFNX1 \ram_reg[119][2]  ( .D(n3118), .CLK(clk), .Q(\ram[119][2] ) );
  DFFNX1 \ram_reg[119][1]  ( .D(n3117), .CLK(clk), .Q(\ram[119][1] ) );
  DFFNX1 \ram_reg[119][0]  ( .D(n3116), .CLK(clk), .Q(\ram[119][0] ) );
  DFFNX1 \ram_reg[120][7]  ( .D(n3115), .CLK(clk), .Q(\ram[120][7] ) );
  DFFNX1 \ram_reg[120][6]  ( .D(n3114), .CLK(clk), .Q(\ram[120][6] ) );
  DFFNX1 \ram_reg[120][5]  ( .D(n3113), .CLK(clk), .Q(\ram[120][5] ) );
  DFFNX1 \ram_reg[120][4]  ( .D(n3112), .CLK(clk), .Q(\ram[120][4] ) );
  DFFNX1 \ram_reg[120][3]  ( .D(n3111), .CLK(clk), .Q(\ram[120][3] ) );
  DFFNX1 \ram_reg[120][2]  ( .D(n3110), .CLK(clk), .Q(\ram[120][2] ) );
  DFFNX1 \ram_reg[120][1]  ( .D(n3109), .CLK(clk), .Q(\ram[120][1] ) );
  DFFNX1 \ram_reg[120][0]  ( .D(n3108), .CLK(clk), .Q(\ram[120][0] ) );
  DFFNX1 \ram_reg[121][7]  ( .D(n3107), .CLK(clk), .Q(\ram[121][7] ) );
  DFFNX1 \ram_reg[121][6]  ( .D(n3106), .CLK(clk), .Q(\ram[121][6] ) );
  DFFNX1 \ram_reg[121][5]  ( .D(n3105), .CLK(clk), .Q(\ram[121][5] ) );
  DFFNX1 \ram_reg[121][4]  ( .D(n3104), .CLK(clk), .Q(\ram[121][4] ) );
  DFFNX1 \ram_reg[121][3]  ( .D(n3103), .CLK(clk), .Q(\ram[121][3] ) );
  DFFNX1 \ram_reg[121][2]  ( .D(n3102), .CLK(clk), .Q(\ram[121][2] ) );
  DFFNX1 \ram_reg[121][1]  ( .D(n3101), .CLK(clk), .Q(\ram[121][1] ) );
  DFFNX1 \ram_reg[121][0]  ( .D(n3100), .CLK(clk), .Q(\ram[121][0] ) );
  DFFNX1 \ram_reg[122][7]  ( .D(n3099), .CLK(clk), .Q(\ram[122][7] ) );
  DFFNX1 \ram_reg[122][6]  ( .D(n3098), .CLK(clk), .Q(\ram[122][6] ) );
  DFFNX1 \ram_reg[122][5]  ( .D(n3097), .CLK(clk), .Q(\ram[122][5] ) );
  DFFNX1 \ram_reg[122][4]  ( .D(n3096), .CLK(clk), .Q(\ram[122][4] ) );
  DFFNX1 \ram_reg[122][3]  ( .D(n3095), .CLK(clk), .Q(\ram[122][3] ) );
  DFFNX1 \ram_reg[122][2]  ( .D(n3094), .CLK(clk), .Q(\ram[122][2] ) );
  DFFNX1 \ram_reg[122][1]  ( .D(n3093), .CLK(clk), .Q(\ram[122][1] ) );
  DFFNX1 \ram_reg[122][0]  ( .D(n3092), .CLK(clk), .Q(\ram[122][0] ) );
  DFFNX1 \ram_reg[123][7]  ( .D(n3091), .CLK(clk), .Q(\ram[123][7] ) );
  DFFNX1 \ram_reg[123][6]  ( .D(n3090), .CLK(clk), .Q(\ram[123][6] ) );
  DFFNX1 \ram_reg[123][5]  ( .D(n3089), .CLK(clk), .Q(\ram[123][5] ) );
  DFFNX1 \ram_reg[123][4]  ( .D(n3088), .CLK(clk), .Q(\ram[123][4] ) );
  DFFNX1 \ram_reg[123][3]  ( .D(n3087), .CLK(clk), .Q(\ram[123][3] ) );
  DFFNX1 \ram_reg[123][2]  ( .D(n3086), .CLK(clk), .Q(\ram[123][2] ) );
  DFFNX1 \ram_reg[123][1]  ( .D(n3085), .CLK(clk), .Q(\ram[123][1] ) );
  DFFNX1 \ram_reg[123][0]  ( .D(n3084), .CLK(clk), .Q(\ram[123][0] ) );
  DFFNX1 \ram_reg[124][7]  ( .D(n3083), .CLK(clk), .Q(\ram[124][7] ) );
  DFFNX1 \ram_reg[124][6]  ( .D(n3082), .CLK(clk), .Q(\ram[124][6] ) );
  DFFNX1 \ram_reg[124][5]  ( .D(n3081), .CLK(clk), .Q(\ram[124][5] ) );
  DFFNX1 \ram_reg[124][4]  ( .D(n3080), .CLK(clk), .Q(\ram[124][4] ) );
  DFFNX1 \ram_reg[124][3]  ( .D(n3079), .CLK(clk), .Q(\ram[124][3] ) );
  DFFNX1 \ram_reg[124][2]  ( .D(n3078), .CLK(clk), .Q(\ram[124][2] ) );
  DFFNX1 \ram_reg[124][1]  ( .D(n3077), .CLK(clk), .Q(\ram[124][1] ) );
  DFFNX1 \ram_reg[124][0]  ( .D(n3076), .CLK(clk), .Q(\ram[124][0] ) );
  DFFNX1 \ram_reg[125][7]  ( .D(n3075), .CLK(clk), .Q(\ram[125][7] ) );
  DFFNX1 \ram_reg[125][6]  ( .D(n3074), .CLK(clk), .Q(\ram[125][6] ) );
  DFFNX1 \ram_reg[125][5]  ( .D(n3073), .CLK(clk), .Q(\ram[125][5] ) );
  DFFNX1 \ram_reg[125][4]  ( .D(n3072), .CLK(clk), .Q(\ram[125][4] ) );
  DFFNX1 \ram_reg[125][3]  ( .D(n3071), .CLK(clk), .Q(\ram[125][3] ) );
  DFFNX1 \ram_reg[125][2]  ( .D(n3070), .CLK(clk), .Q(\ram[125][2] ) );
  DFFNX1 \ram_reg[125][1]  ( .D(n3069), .CLK(clk), .Q(\ram[125][1] ) );
  DFFNX1 \ram_reg[125][0]  ( .D(n3068), .CLK(clk), .Q(\ram[125][0] ) );
  DFFNX1 \ram_reg[126][7]  ( .D(n3067), .CLK(clk), .Q(\ram[126][7] ) );
  DFFNX1 \ram_reg[126][6]  ( .D(n3066), .CLK(clk), .Q(\ram[126][6] ) );
  DFFNX1 \ram_reg[126][5]  ( .D(n3065), .CLK(clk), .Q(\ram[126][5] ) );
  DFFNX1 \ram_reg[126][4]  ( .D(n3064), .CLK(clk), .Q(\ram[126][4] ) );
  DFFNX1 \ram_reg[126][3]  ( .D(n3063), .CLK(clk), .Q(\ram[126][3] ) );
  DFFNX1 \ram_reg[126][2]  ( .D(n3062), .CLK(clk), .Q(\ram[126][2] ) );
  DFFNX1 \ram_reg[126][1]  ( .D(n3061), .CLK(clk), .Q(\ram[126][1] ) );
  DFFNX1 \ram_reg[126][0]  ( .D(n3060), .CLK(clk), .Q(\ram[126][0] ) );
  DFFNX1 \ram_reg[127][7]  ( .D(n3059), .CLK(clk), .Q(\ram[127][7] ) );
  DFFNX1 \ram_reg[127][6]  ( .D(n3058), .CLK(clk), .Q(\ram[127][6] ) );
  DFFNX1 \ram_reg[127][5]  ( .D(n3057), .CLK(clk), .Q(\ram[127][5] ) );
  DFFNX1 \ram_reg[127][4]  ( .D(n3056), .CLK(clk), .Q(\ram[127][4] ) );
  DFFNX1 \ram_reg[127][3]  ( .D(n3055), .CLK(clk), .Q(\ram[127][3] ) );
  DFFNX1 \ram_reg[127][2]  ( .D(n3054), .CLK(clk), .Q(\ram[127][2] ) );
  DFFNX1 \ram_reg[127][1]  ( .D(n3053), .CLK(clk), .Q(\ram[127][1] ) );
  DFFNX1 \ram_reg[127][0]  ( .D(n3052), .CLK(clk), .Q(\ram[127][0] ) );
  DFFNX1 \ram_reg[128][7]  ( .D(n3051), .CLK(clk), .Q(\ram[128][7] ) );
  DFFNX1 \ram_reg[128][6]  ( .D(n3050), .CLK(clk), .Q(\ram[128][6] ) );
  DFFNX1 \ram_reg[128][5]  ( .D(n3049), .CLK(clk), .Q(\ram[128][5] ) );
  DFFNX1 \ram_reg[128][4]  ( .D(n3048), .CLK(clk), .Q(\ram[128][4] ) );
  DFFNX1 \ram_reg[128][3]  ( .D(n3047), .CLK(clk), .Q(\ram[128][3] ) );
  DFFNX1 \ram_reg[128][2]  ( .D(n3046), .CLK(clk), .Q(\ram[128][2] ) );
  DFFNX1 \ram_reg[128][1]  ( .D(n3045), .CLK(clk), .Q(\ram[128][1] ) );
  DFFNX1 \ram_reg[128][0]  ( .D(n3044), .CLK(clk), .Q(\ram[128][0] ) );
  DFFNX1 \ram_reg[129][7]  ( .D(n3043), .CLK(clk), .Q(\ram[129][7] ) );
  DFFNX1 \ram_reg[129][6]  ( .D(n3042), .CLK(clk), .Q(\ram[129][6] ) );
  DFFNX1 \ram_reg[129][5]  ( .D(n3041), .CLK(clk), .Q(\ram[129][5] ) );
  DFFNX1 \ram_reg[129][4]  ( .D(n3040), .CLK(clk), .Q(\ram[129][4] ) );
  DFFNX1 \ram_reg[129][3]  ( .D(n3039), .CLK(clk), .Q(\ram[129][3] ) );
  DFFNX1 \ram_reg[129][2]  ( .D(n3038), .CLK(clk), .Q(\ram[129][2] ) );
  DFFNX1 \ram_reg[129][1]  ( .D(n3037), .CLK(clk), .Q(\ram[129][1] ) );
  DFFNX1 \ram_reg[129][0]  ( .D(n3036), .CLK(clk), .Q(\ram[129][0] ) );
  DFFNX1 \ram_reg[130][7]  ( .D(n3035), .CLK(clk), .Q(\ram[130][7] ) );
  DFFNX1 \ram_reg[130][6]  ( .D(n3034), .CLK(clk), .Q(\ram[130][6] ) );
  DFFNX1 \ram_reg[130][5]  ( .D(n3033), .CLK(clk), .Q(\ram[130][5] ) );
  DFFNX1 \ram_reg[130][4]  ( .D(n3032), .CLK(clk), .Q(\ram[130][4] ) );
  DFFNX1 \ram_reg[130][3]  ( .D(n3031), .CLK(clk), .Q(\ram[130][3] ) );
  DFFNX1 \ram_reg[130][2]  ( .D(n3030), .CLK(clk), .Q(\ram[130][2] ) );
  DFFNX1 \ram_reg[130][1]  ( .D(n3029), .CLK(clk), .Q(\ram[130][1] ) );
  DFFNX1 \ram_reg[130][0]  ( .D(n3028), .CLK(clk), .Q(\ram[130][0] ) );
  DFFNX1 \ram_reg[131][7]  ( .D(n3027), .CLK(clk), .Q(\ram[131][7] ) );
  DFFNX1 \ram_reg[131][6]  ( .D(n3026), .CLK(clk), .Q(\ram[131][6] ) );
  DFFNX1 \ram_reg[131][5]  ( .D(n3025), .CLK(clk), .Q(\ram[131][5] ) );
  DFFNX1 \ram_reg[131][4]  ( .D(n3024), .CLK(clk), .Q(\ram[131][4] ) );
  DFFNX1 \ram_reg[131][3]  ( .D(n3023), .CLK(clk), .Q(\ram[131][3] ) );
  DFFNX1 \ram_reg[131][2]  ( .D(n3022), .CLK(clk), .Q(\ram[131][2] ) );
  DFFNX1 \ram_reg[131][1]  ( .D(n3021), .CLK(clk), .Q(\ram[131][1] ) );
  DFFNX1 \ram_reg[131][0]  ( .D(n3020), .CLK(clk), .Q(\ram[131][0] ) );
  DFFNX1 \ram_reg[132][7]  ( .D(n3019), .CLK(clk), .Q(\ram[132][7] ) );
  DFFNX1 \ram_reg[132][6]  ( .D(n3018), .CLK(clk), .Q(\ram[132][6] ) );
  DFFNX1 \ram_reg[132][5]  ( .D(n3017), .CLK(clk), .Q(\ram[132][5] ) );
  DFFNX1 \ram_reg[132][4]  ( .D(n3016), .CLK(clk), .Q(\ram[132][4] ) );
  DFFNX1 \ram_reg[132][3]  ( .D(n3015), .CLK(clk), .Q(\ram[132][3] ) );
  DFFNX1 \ram_reg[132][2]  ( .D(n3014), .CLK(clk), .Q(\ram[132][2] ) );
  DFFNX1 \ram_reg[132][1]  ( .D(n3013), .CLK(clk), .Q(\ram[132][1] ) );
  DFFNX1 \ram_reg[132][0]  ( .D(n3012), .CLK(clk), .Q(\ram[132][0] ) );
  DFFNX1 \ram_reg[133][7]  ( .D(n3011), .CLK(clk), .Q(\ram[133][7] ) );
  DFFNX1 \ram_reg[133][6]  ( .D(n3010), .CLK(clk), .Q(\ram[133][6] ) );
  DFFNX1 \ram_reg[133][5]  ( .D(n3009), .CLK(clk), .Q(\ram[133][5] ) );
  DFFNX1 \ram_reg[133][4]  ( .D(n3008), .CLK(clk), .Q(\ram[133][4] ) );
  DFFNX1 \ram_reg[133][3]  ( .D(n3007), .CLK(clk), .Q(\ram[133][3] ) );
  DFFNX1 \ram_reg[133][2]  ( .D(n3006), .CLK(clk), .Q(\ram[133][2] ) );
  DFFNX1 \ram_reg[133][1]  ( .D(n3005), .CLK(clk), .Q(\ram[133][1] ) );
  DFFNX1 \ram_reg[133][0]  ( .D(n3004), .CLK(clk), .Q(\ram[133][0] ) );
  DFFNX1 \ram_reg[134][7]  ( .D(n3003), .CLK(clk), .Q(\ram[134][7] ) );
  DFFNX1 \ram_reg[134][6]  ( .D(n3002), .CLK(clk), .Q(\ram[134][6] ) );
  DFFNX1 \ram_reg[134][5]  ( .D(n3001), .CLK(clk), .Q(\ram[134][5] ) );
  DFFNX1 \ram_reg[134][4]  ( .D(n3000), .CLK(clk), .Q(\ram[134][4] ) );
  DFFNX1 \ram_reg[134][3]  ( .D(n2999), .CLK(clk), .Q(\ram[134][3] ) );
  DFFNX1 \ram_reg[134][2]  ( .D(n2998), .CLK(clk), .Q(\ram[134][2] ) );
  DFFNX1 \ram_reg[134][1]  ( .D(n2997), .CLK(clk), .Q(\ram[134][1] ) );
  DFFNX1 \ram_reg[134][0]  ( .D(n2996), .CLK(clk), .Q(\ram[134][0] ) );
  DFFNX1 \ram_reg[135][7]  ( .D(n2995), .CLK(clk), .Q(\ram[135][7] ) );
  DFFNX1 \ram_reg[135][6]  ( .D(n2994), .CLK(clk), .Q(\ram[135][6] ) );
  DFFNX1 \ram_reg[135][5]  ( .D(n2993), .CLK(clk), .Q(\ram[135][5] ) );
  DFFNX1 \ram_reg[135][4]  ( .D(n2992), .CLK(clk), .Q(\ram[135][4] ) );
  DFFNX1 \ram_reg[135][3]  ( .D(n2991), .CLK(clk), .Q(\ram[135][3] ) );
  DFFNX1 \ram_reg[135][2]  ( .D(n2990), .CLK(clk), .Q(\ram[135][2] ) );
  DFFNX1 \ram_reg[135][1]  ( .D(n2989), .CLK(clk), .Q(\ram[135][1] ) );
  DFFNX1 \ram_reg[135][0]  ( .D(n2988), .CLK(clk), .Q(\ram[135][0] ) );
  DFFNX1 \ram_reg[136][7]  ( .D(n2987), .CLK(clk), .Q(\ram[136][7] ) );
  DFFNX1 \ram_reg[136][6]  ( .D(n2986), .CLK(clk), .Q(\ram[136][6] ) );
  DFFNX1 \ram_reg[136][5]  ( .D(n2985), .CLK(clk), .Q(\ram[136][5] ) );
  DFFNX1 \ram_reg[136][4]  ( .D(n2984), .CLK(clk), .Q(\ram[136][4] ) );
  DFFNX1 \ram_reg[136][3]  ( .D(n2983), .CLK(clk), .Q(\ram[136][3] ) );
  DFFNX1 \ram_reg[136][2]  ( .D(n2982), .CLK(clk), .Q(\ram[136][2] ) );
  DFFNX1 \ram_reg[136][1]  ( .D(n2981), .CLK(clk), .Q(\ram[136][1] ) );
  DFFNX1 \ram_reg[136][0]  ( .D(n2980), .CLK(clk), .Q(\ram[136][0] ) );
  DFFNX1 \ram_reg[137][7]  ( .D(n2979), .CLK(clk), .Q(\ram[137][7] ) );
  DFFNX1 \ram_reg[137][6]  ( .D(n2978), .CLK(clk), .Q(\ram[137][6] ) );
  DFFNX1 \ram_reg[137][5]  ( .D(n2977), .CLK(clk), .Q(\ram[137][5] ) );
  DFFNX1 \ram_reg[137][4]  ( .D(n2976), .CLK(clk), .Q(\ram[137][4] ) );
  DFFNX1 \ram_reg[137][3]  ( .D(n2975), .CLK(clk), .Q(\ram[137][3] ) );
  DFFNX1 \ram_reg[137][2]  ( .D(n2974), .CLK(clk), .Q(\ram[137][2] ) );
  DFFNX1 \ram_reg[137][1]  ( .D(n2973), .CLK(clk), .Q(\ram[137][1] ) );
  DFFNX1 \ram_reg[137][0]  ( .D(n2972), .CLK(clk), .Q(\ram[137][0] ) );
  DFFNX1 \ram_reg[138][7]  ( .D(n2971), .CLK(clk), .Q(\ram[138][7] ) );
  DFFNX1 \ram_reg[138][6]  ( .D(n2970), .CLK(clk), .Q(\ram[138][6] ) );
  DFFNX1 \ram_reg[138][5]  ( .D(n2969), .CLK(clk), .Q(\ram[138][5] ) );
  DFFNX1 \ram_reg[138][4]  ( .D(n2968), .CLK(clk), .Q(\ram[138][4] ) );
  DFFNX1 \ram_reg[138][3]  ( .D(n2967), .CLK(clk), .Q(\ram[138][3] ) );
  DFFNX1 \ram_reg[138][2]  ( .D(n2966), .CLK(clk), .Q(\ram[138][2] ) );
  DFFNX1 \ram_reg[138][1]  ( .D(n2965), .CLK(clk), .Q(\ram[138][1] ) );
  DFFNX1 \ram_reg[138][0]  ( .D(n2964), .CLK(clk), .Q(\ram[138][0] ) );
  DFFNX1 \ram_reg[139][7]  ( .D(n2963), .CLK(clk), .Q(\ram[139][7] ) );
  DFFNX1 \ram_reg[139][6]  ( .D(n2962), .CLK(clk), .Q(\ram[139][6] ) );
  DFFNX1 \ram_reg[139][5]  ( .D(n2961), .CLK(clk), .Q(\ram[139][5] ) );
  DFFNX1 \ram_reg[139][4]  ( .D(n2960), .CLK(clk), .Q(\ram[139][4] ) );
  DFFNX1 \ram_reg[139][3]  ( .D(n2959), .CLK(clk), .Q(\ram[139][3] ) );
  DFFNX1 \ram_reg[139][2]  ( .D(n2958), .CLK(clk), .Q(\ram[139][2] ) );
  DFFNX1 \ram_reg[139][1]  ( .D(n2957), .CLK(clk), .Q(\ram[139][1] ) );
  DFFNX1 \ram_reg[139][0]  ( .D(n2956), .CLK(clk), .Q(\ram[139][0] ) );
  DFFNX1 \ram_reg[140][7]  ( .D(n2955), .CLK(clk), .Q(\ram[140][7] ) );
  DFFNX1 \ram_reg[140][6]  ( .D(n2954), .CLK(clk), .Q(\ram[140][6] ) );
  DFFNX1 \ram_reg[140][5]  ( .D(n2953), .CLK(clk), .Q(\ram[140][5] ) );
  DFFNX1 \ram_reg[140][4]  ( .D(n2952), .CLK(clk), .Q(\ram[140][4] ) );
  DFFNX1 \ram_reg[140][3]  ( .D(n2951), .CLK(clk), .Q(\ram[140][3] ) );
  DFFNX1 \ram_reg[140][2]  ( .D(n2950), .CLK(clk), .Q(\ram[140][2] ) );
  DFFNX1 \ram_reg[140][1]  ( .D(n2949), .CLK(clk), .Q(\ram[140][1] ) );
  DFFNX1 \ram_reg[140][0]  ( .D(n2948), .CLK(clk), .Q(\ram[140][0] ) );
  DFFNX1 \ram_reg[141][7]  ( .D(n2947), .CLK(clk), .Q(\ram[141][7] ) );
  DFFNX1 \ram_reg[141][6]  ( .D(n2946), .CLK(clk), .Q(\ram[141][6] ) );
  DFFNX1 \ram_reg[141][5]  ( .D(n2945), .CLK(clk), .Q(\ram[141][5] ) );
  DFFNX1 \ram_reg[141][4]  ( .D(n2944), .CLK(clk), .Q(\ram[141][4] ) );
  DFFNX1 \ram_reg[141][3]  ( .D(n2943), .CLK(clk), .Q(\ram[141][3] ) );
  DFFNX1 \ram_reg[141][2]  ( .D(n2942), .CLK(clk), .Q(\ram[141][2] ) );
  DFFNX1 \ram_reg[141][1]  ( .D(n2941), .CLK(clk), .Q(\ram[141][1] ) );
  DFFNX1 \ram_reg[141][0]  ( .D(n2940), .CLK(clk), .Q(\ram[141][0] ) );
  DFFNX1 \ram_reg[142][7]  ( .D(n2939), .CLK(clk), .Q(\ram[142][7] ) );
  DFFNX1 \ram_reg[142][6]  ( .D(n2938), .CLK(clk), .Q(\ram[142][6] ) );
  DFFNX1 \ram_reg[142][5]  ( .D(n2937), .CLK(clk), .Q(\ram[142][5] ) );
  DFFNX1 \ram_reg[142][4]  ( .D(n2936), .CLK(clk), .Q(\ram[142][4] ) );
  DFFNX1 \ram_reg[142][3]  ( .D(n2935), .CLK(clk), .Q(\ram[142][3] ) );
  DFFNX1 \ram_reg[142][2]  ( .D(n2934), .CLK(clk), .Q(\ram[142][2] ) );
  DFFNX1 \ram_reg[142][1]  ( .D(n2933), .CLK(clk), .Q(\ram[142][1] ) );
  DFFNX1 \ram_reg[142][0]  ( .D(n2932), .CLK(clk), .Q(\ram[142][0] ) );
  DFFNX1 \ram_reg[143][7]  ( .D(n2931), .CLK(clk), .Q(\ram[143][7] ) );
  DFFNX1 \ram_reg[143][6]  ( .D(n2930), .CLK(clk), .Q(\ram[143][6] ) );
  DFFNX1 \ram_reg[143][5]  ( .D(n2929), .CLK(clk), .Q(\ram[143][5] ) );
  DFFNX1 \ram_reg[143][4]  ( .D(n2928), .CLK(clk), .Q(\ram[143][4] ) );
  DFFNX1 \ram_reg[143][3]  ( .D(n2927), .CLK(clk), .Q(\ram[143][3] ) );
  DFFNX1 \ram_reg[143][2]  ( .D(n2926), .CLK(clk), .Q(\ram[143][2] ) );
  DFFNX1 \ram_reg[143][1]  ( .D(n2925), .CLK(clk), .Q(\ram[143][1] ) );
  DFFNX1 \ram_reg[143][0]  ( .D(n2924), .CLK(clk), .Q(\ram[143][0] ) );
  DFFNX1 \ram_reg[144][7]  ( .D(n2923), .CLK(clk), .Q(\ram[144][7] ) );
  DFFNX1 \ram_reg[144][6]  ( .D(n2922), .CLK(clk), .Q(\ram[144][6] ) );
  DFFNX1 \ram_reg[144][5]  ( .D(n2921), .CLK(clk), .Q(\ram[144][5] ) );
  DFFNX1 \ram_reg[144][4]  ( .D(n2920), .CLK(clk), .Q(\ram[144][4] ) );
  DFFNX1 \ram_reg[144][3]  ( .D(n2919), .CLK(clk), .Q(\ram[144][3] ) );
  DFFNX1 \ram_reg[144][2]  ( .D(n2918), .CLK(clk), .Q(\ram[144][2] ) );
  DFFNX1 \ram_reg[144][1]  ( .D(n2917), .CLK(clk), .Q(\ram[144][1] ) );
  DFFNX1 \ram_reg[144][0]  ( .D(n2916), .CLK(clk), .Q(\ram[144][0] ) );
  DFFNX1 \ram_reg[145][7]  ( .D(n2915), .CLK(clk), .Q(\ram[145][7] ) );
  DFFNX1 \ram_reg[145][6]  ( .D(n2914), .CLK(clk), .Q(\ram[145][6] ) );
  DFFNX1 \ram_reg[145][5]  ( .D(n2913), .CLK(clk), .Q(\ram[145][5] ) );
  DFFNX1 \ram_reg[145][4]  ( .D(n2912), .CLK(clk), .Q(\ram[145][4] ) );
  DFFNX1 \ram_reg[145][3]  ( .D(n2911), .CLK(clk), .Q(\ram[145][3] ) );
  DFFNX1 \ram_reg[145][2]  ( .D(n2910), .CLK(clk), .Q(\ram[145][2] ) );
  DFFNX1 \ram_reg[145][1]  ( .D(n2909), .CLK(clk), .Q(\ram[145][1] ) );
  DFFNX1 \ram_reg[145][0]  ( .D(n2908), .CLK(clk), .Q(\ram[145][0] ) );
  DFFNX1 \ram_reg[146][7]  ( .D(n2907), .CLK(clk), .Q(\ram[146][7] ) );
  DFFNX1 \ram_reg[146][6]  ( .D(n2906), .CLK(clk), .Q(\ram[146][6] ) );
  DFFNX1 \ram_reg[146][5]  ( .D(n2905), .CLK(clk), .Q(\ram[146][5] ) );
  DFFNX1 \ram_reg[146][4]  ( .D(n2904), .CLK(clk), .Q(\ram[146][4] ) );
  DFFNX1 \ram_reg[146][3]  ( .D(n2903), .CLK(clk), .Q(\ram[146][3] ) );
  DFFNX1 \ram_reg[146][2]  ( .D(n2902), .CLK(clk), .Q(\ram[146][2] ) );
  DFFNX1 \ram_reg[146][1]  ( .D(n2901), .CLK(clk), .Q(\ram[146][1] ) );
  DFFNX1 \ram_reg[146][0]  ( .D(n2900), .CLK(clk), .Q(\ram[146][0] ) );
  DFFNX1 \ram_reg[147][7]  ( .D(n2899), .CLK(clk), .Q(\ram[147][7] ) );
  DFFNX1 \ram_reg[147][6]  ( .D(n2898), .CLK(clk), .Q(\ram[147][6] ) );
  DFFNX1 \ram_reg[147][5]  ( .D(n2897), .CLK(clk), .Q(\ram[147][5] ) );
  DFFNX1 \ram_reg[147][4]  ( .D(n2896), .CLK(clk), .Q(\ram[147][4] ) );
  DFFNX1 \ram_reg[147][3]  ( .D(n2895), .CLK(clk), .Q(\ram[147][3] ) );
  DFFNX1 \ram_reg[147][2]  ( .D(n2894), .CLK(clk), .Q(\ram[147][2] ) );
  DFFNX1 \ram_reg[147][1]  ( .D(n2893), .CLK(clk), .Q(\ram[147][1] ) );
  DFFNX1 \ram_reg[147][0]  ( .D(n2892), .CLK(clk), .Q(\ram[147][0] ) );
  DFFNX1 \ram_reg[148][7]  ( .D(n2891), .CLK(clk), .Q(\ram[148][7] ) );
  DFFNX1 \ram_reg[148][6]  ( .D(n2890), .CLK(clk), .Q(\ram[148][6] ) );
  DFFNX1 \ram_reg[148][5]  ( .D(n2889), .CLK(clk), .Q(\ram[148][5] ) );
  DFFNX1 \ram_reg[148][4]  ( .D(n2888), .CLK(clk), .Q(\ram[148][4] ) );
  DFFNX1 \ram_reg[148][3]  ( .D(n2887), .CLK(clk), .Q(\ram[148][3] ) );
  DFFNX1 \ram_reg[148][2]  ( .D(n2886), .CLK(clk), .Q(\ram[148][2] ) );
  DFFNX1 \ram_reg[148][1]  ( .D(n2885), .CLK(clk), .Q(\ram[148][1] ) );
  DFFNX1 \ram_reg[148][0]  ( .D(n2884), .CLK(clk), .Q(\ram[148][0] ) );
  DFFNX1 \ram_reg[149][7]  ( .D(n2883), .CLK(clk), .Q(\ram[149][7] ) );
  DFFNX1 \ram_reg[149][6]  ( .D(n2882), .CLK(clk), .Q(\ram[149][6] ) );
  DFFNX1 \ram_reg[149][5]  ( .D(n2881), .CLK(clk), .Q(\ram[149][5] ) );
  DFFNX1 \ram_reg[149][4]  ( .D(n2880), .CLK(clk), .Q(\ram[149][4] ) );
  DFFNX1 \ram_reg[149][3]  ( .D(n2879), .CLK(clk), .Q(\ram[149][3] ) );
  DFFNX1 \ram_reg[149][2]  ( .D(n2878), .CLK(clk), .Q(\ram[149][2] ) );
  DFFNX1 \ram_reg[149][1]  ( .D(n2877), .CLK(clk), .Q(\ram[149][1] ) );
  DFFNX1 \ram_reg[149][0]  ( .D(n2876), .CLK(clk), .Q(\ram[149][0] ) );
  DFFNX1 \ram_reg[150][7]  ( .D(n2875), .CLK(clk), .Q(\ram[150][7] ) );
  DFFNX1 \ram_reg[150][6]  ( .D(n2874), .CLK(clk), .Q(\ram[150][6] ) );
  DFFNX1 \ram_reg[150][5]  ( .D(n2873), .CLK(clk), .Q(\ram[150][5] ) );
  DFFNX1 \ram_reg[150][4]  ( .D(n2872), .CLK(clk), .Q(\ram[150][4] ) );
  DFFNX1 \ram_reg[150][3]  ( .D(n2871), .CLK(clk), .Q(\ram[150][3] ) );
  DFFNX1 \ram_reg[150][2]  ( .D(n2870), .CLK(clk), .Q(\ram[150][2] ) );
  DFFNX1 \ram_reg[150][1]  ( .D(n2869), .CLK(clk), .Q(\ram[150][1] ) );
  DFFNX1 \ram_reg[150][0]  ( .D(n2868), .CLK(clk), .Q(\ram[150][0] ) );
  DFFNX1 \ram_reg[151][7]  ( .D(n2867), .CLK(clk), .Q(\ram[151][7] ) );
  DFFNX1 \ram_reg[151][6]  ( .D(n2866), .CLK(clk), .Q(\ram[151][6] ) );
  DFFNX1 \ram_reg[151][5]  ( .D(n2865), .CLK(clk), .Q(\ram[151][5] ) );
  DFFNX1 \ram_reg[151][4]  ( .D(n2864), .CLK(clk), .Q(\ram[151][4] ) );
  DFFNX1 \ram_reg[151][3]  ( .D(n2863), .CLK(clk), .Q(\ram[151][3] ) );
  DFFNX1 \ram_reg[151][2]  ( .D(n2862), .CLK(clk), .Q(\ram[151][2] ) );
  DFFNX1 \ram_reg[151][1]  ( .D(n2861), .CLK(clk), .Q(\ram[151][1] ) );
  DFFNX1 \ram_reg[151][0]  ( .D(n2860), .CLK(clk), .Q(\ram[151][0] ) );
  DFFNX1 \ram_reg[152][7]  ( .D(n2859), .CLK(clk), .Q(\ram[152][7] ) );
  DFFNX1 \ram_reg[152][6]  ( .D(n2858), .CLK(clk), .Q(\ram[152][6] ) );
  DFFNX1 \ram_reg[152][5]  ( .D(n2857), .CLK(clk), .Q(\ram[152][5] ) );
  DFFNX1 \ram_reg[152][4]  ( .D(n2856), .CLK(clk), .Q(\ram[152][4] ) );
  DFFNX1 \ram_reg[152][3]  ( .D(n2855), .CLK(clk), .Q(\ram[152][3] ) );
  DFFNX1 \ram_reg[152][2]  ( .D(n2854), .CLK(clk), .Q(\ram[152][2] ) );
  DFFNX1 \ram_reg[152][1]  ( .D(n2853), .CLK(clk), .Q(\ram[152][1] ) );
  DFFNX1 \ram_reg[152][0]  ( .D(n2852), .CLK(clk), .Q(\ram[152][0] ) );
  DFFNX1 \ram_reg[153][7]  ( .D(n2851), .CLK(clk), .Q(\ram[153][7] ) );
  DFFNX1 \ram_reg[153][6]  ( .D(n2850), .CLK(clk), .Q(\ram[153][6] ) );
  DFFNX1 \ram_reg[153][5]  ( .D(n2849), .CLK(clk), .Q(\ram[153][5] ) );
  DFFNX1 \ram_reg[153][4]  ( .D(n2848), .CLK(clk), .Q(\ram[153][4] ) );
  DFFNX1 \ram_reg[153][3]  ( .D(n2847), .CLK(clk), .Q(\ram[153][3] ) );
  DFFNX1 \ram_reg[153][2]  ( .D(n2846), .CLK(clk), .Q(\ram[153][2] ) );
  DFFNX1 \ram_reg[153][1]  ( .D(n2845), .CLK(clk), .Q(\ram[153][1] ) );
  DFFNX1 \ram_reg[153][0]  ( .D(n2844), .CLK(clk), .Q(\ram[153][0] ) );
  DFFNX1 \ram_reg[154][7]  ( .D(n2843), .CLK(clk), .Q(\ram[154][7] ) );
  DFFNX1 \ram_reg[154][6]  ( .D(n2842), .CLK(clk), .Q(\ram[154][6] ) );
  DFFNX1 \ram_reg[154][5]  ( .D(n2841), .CLK(clk), .Q(\ram[154][5] ) );
  DFFNX1 \ram_reg[154][4]  ( .D(n2840), .CLK(clk), .Q(\ram[154][4] ) );
  DFFNX1 \ram_reg[154][3]  ( .D(n2839), .CLK(clk), .Q(\ram[154][3] ) );
  DFFNX1 \ram_reg[154][2]  ( .D(n2838), .CLK(clk), .Q(\ram[154][2] ) );
  DFFNX1 \ram_reg[154][1]  ( .D(n2837), .CLK(clk), .Q(\ram[154][1] ) );
  DFFNX1 \ram_reg[154][0]  ( .D(n2836), .CLK(clk), .Q(\ram[154][0] ) );
  DFFNX1 \ram_reg[155][7]  ( .D(n2835), .CLK(clk), .Q(\ram[155][7] ) );
  DFFNX1 \ram_reg[155][6]  ( .D(n2834), .CLK(clk), .Q(\ram[155][6] ) );
  DFFNX1 \ram_reg[155][5]  ( .D(n2833), .CLK(clk), .Q(\ram[155][5] ) );
  DFFNX1 \ram_reg[155][4]  ( .D(n2832), .CLK(clk), .Q(\ram[155][4] ) );
  DFFNX1 \ram_reg[155][3]  ( .D(n2831), .CLK(clk), .Q(\ram[155][3] ) );
  DFFNX1 \ram_reg[155][2]  ( .D(n2830), .CLK(clk), .Q(\ram[155][2] ) );
  DFFNX1 \ram_reg[155][1]  ( .D(n2829), .CLK(clk), .Q(\ram[155][1] ) );
  DFFNX1 \ram_reg[155][0]  ( .D(n2828), .CLK(clk), .Q(\ram[155][0] ) );
  DFFNX1 \ram_reg[156][7]  ( .D(n2827), .CLK(clk), .Q(\ram[156][7] ) );
  DFFNX1 \ram_reg[156][6]  ( .D(n2826), .CLK(clk), .Q(\ram[156][6] ) );
  DFFNX1 \ram_reg[156][5]  ( .D(n2825), .CLK(clk), .Q(\ram[156][5] ) );
  DFFNX1 \ram_reg[156][4]  ( .D(n2824), .CLK(clk), .Q(\ram[156][4] ) );
  DFFNX1 \ram_reg[156][3]  ( .D(n2823), .CLK(clk), .Q(\ram[156][3] ) );
  DFFNX1 \ram_reg[156][2]  ( .D(n2822), .CLK(clk), .Q(\ram[156][2] ) );
  DFFNX1 \ram_reg[156][1]  ( .D(n2821), .CLK(clk), .Q(\ram[156][1] ) );
  DFFNX1 \ram_reg[156][0]  ( .D(n2820), .CLK(clk), .Q(\ram[156][0] ) );
  DFFNX1 \ram_reg[157][7]  ( .D(n2819), .CLK(clk), .Q(\ram[157][7] ) );
  DFFNX1 \ram_reg[157][6]  ( .D(n2818), .CLK(clk), .Q(\ram[157][6] ) );
  DFFNX1 \ram_reg[157][5]  ( .D(n2817), .CLK(clk), .Q(\ram[157][5] ) );
  DFFNX1 \ram_reg[157][4]  ( .D(n2816), .CLK(clk), .Q(\ram[157][4] ) );
  DFFNX1 \ram_reg[157][3]  ( .D(n2815), .CLK(clk), .Q(\ram[157][3] ) );
  DFFNX1 \ram_reg[157][2]  ( .D(n2814), .CLK(clk), .Q(\ram[157][2] ) );
  DFFNX1 \ram_reg[157][1]  ( .D(n2813), .CLK(clk), .Q(\ram[157][1] ) );
  DFFNX1 \ram_reg[157][0]  ( .D(n2812), .CLK(clk), .Q(\ram[157][0] ) );
  DFFNX1 \ram_reg[158][7]  ( .D(n2811), .CLK(clk), .Q(\ram[158][7] ) );
  DFFNX1 \ram_reg[158][6]  ( .D(n2810), .CLK(clk), .Q(\ram[158][6] ) );
  DFFNX1 \ram_reg[158][5]  ( .D(n2809), .CLK(clk), .Q(\ram[158][5] ) );
  DFFNX1 \ram_reg[158][4]  ( .D(n2808), .CLK(clk), .Q(\ram[158][4] ) );
  DFFNX1 \ram_reg[158][3]  ( .D(n2807), .CLK(clk), .Q(\ram[158][3] ) );
  DFFNX1 \ram_reg[158][2]  ( .D(n2806), .CLK(clk), .Q(\ram[158][2] ) );
  DFFNX1 \ram_reg[158][1]  ( .D(n2805), .CLK(clk), .Q(\ram[158][1] ) );
  DFFNX1 \ram_reg[158][0]  ( .D(n2804), .CLK(clk), .Q(\ram[158][0] ) );
  DFFNX1 \ram_reg[159][7]  ( .D(n2803), .CLK(clk), .Q(\ram[159][7] ) );
  DFFNX1 \ram_reg[159][6]  ( .D(n2802), .CLK(clk), .Q(\ram[159][6] ) );
  DFFNX1 \ram_reg[159][5]  ( .D(n2801), .CLK(clk), .Q(\ram[159][5] ) );
  DFFNX1 \ram_reg[159][4]  ( .D(n2800), .CLK(clk), .Q(\ram[159][4] ) );
  DFFNX1 \ram_reg[159][3]  ( .D(n2799), .CLK(clk), .Q(\ram[159][3] ) );
  DFFNX1 \ram_reg[159][2]  ( .D(n2798), .CLK(clk), .Q(\ram[159][2] ) );
  DFFNX1 \ram_reg[159][1]  ( .D(n2797), .CLK(clk), .Q(\ram[159][1] ) );
  DFFNX1 \ram_reg[159][0]  ( .D(n2796), .CLK(clk), .Q(\ram[159][0] ) );
  DFFNX1 \ram_reg[160][7]  ( .D(n2795), .CLK(clk), .Q(\ram[160][7] ) );
  DFFNX1 \ram_reg[160][6]  ( .D(n2794), .CLK(clk), .Q(\ram[160][6] ) );
  DFFNX1 \ram_reg[160][5]  ( .D(n2793), .CLK(clk), .Q(\ram[160][5] ) );
  DFFNX1 \ram_reg[160][4]  ( .D(n2792), .CLK(clk), .Q(\ram[160][4] ) );
  DFFNX1 \ram_reg[160][3]  ( .D(n2791), .CLK(clk), .Q(\ram[160][3] ) );
  DFFNX1 \ram_reg[160][2]  ( .D(n2790), .CLK(clk), .Q(\ram[160][2] ) );
  DFFNX1 \ram_reg[160][1]  ( .D(n2789), .CLK(clk), .Q(\ram[160][1] ) );
  DFFNX1 \ram_reg[160][0]  ( .D(n2788), .CLK(clk), .Q(\ram[160][0] ) );
  DFFNX1 \ram_reg[161][7]  ( .D(n2787), .CLK(clk), .Q(\ram[161][7] ) );
  DFFNX1 \ram_reg[161][6]  ( .D(n2786), .CLK(clk), .Q(\ram[161][6] ) );
  DFFNX1 \ram_reg[161][5]  ( .D(n2785), .CLK(clk), .Q(\ram[161][5] ) );
  DFFNX1 \ram_reg[161][4]  ( .D(n2784), .CLK(clk), .Q(\ram[161][4] ) );
  DFFNX1 \ram_reg[161][3]  ( .D(n2783), .CLK(clk), .Q(\ram[161][3] ) );
  DFFNX1 \ram_reg[161][2]  ( .D(n2782), .CLK(clk), .Q(\ram[161][2] ) );
  DFFNX1 \ram_reg[161][1]  ( .D(n2781), .CLK(clk), .Q(\ram[161][1] ) );
  DFFNX1 \ram_reg[161][0]  ( .D(n2780), .CLK(clk), .Q(\ram[161][0] ) );
  DFFNX1 \ram_reg[162][7]  ( .D(n2779), .CLK(clk), .Q(\ram[162][7] ) );
  DFFNX1 \ram_reg[162][6]  ( .D(n2778), .CLK(clk), .Q(\ram[162][6] ) );
  DFFNX1 \ram_reg[162][5]  ( .D(n2777), .CLK(clk), .Q(\ram[162][5] ) );
  DFFNX1 \ram_reg[162][4]  ( .D(n2776), .CLK(clk), .Q(\ram[162][4] ) );
  DFFNX1 \ram_reg[162][3]  ( .D(n2775), .CLK(clk), .Q(\ram[162][3] ) );
  DFFNX1 \ram_reg[162][2]  ( .D(n2774), .CLK(clk), .Q(\ram[162][2] ) );
  DFFNX1 \ram_reg[162][1]  ( .D(n2773), .CLK(clk), .Q(\ram[162][1] ) );
  DFFNX1 \ram_reg[162][0]  ( .D(n2772), .CLK(clk), .Q(\ram[162][0] ) );
  DFFNX1 \ram_reg[163][7]  ( .D(n2771), .CLK(clk), .Q(\ram[163][7] ) );
  DFFNX1 \ram_reg[163][6]  ( .D(n2770), .CLK(clk), .Q(\ram[163][6] ) );
  DFFNX1 \ram_reg[163][5]  ( .D(n2769), .CLK(clk), .Q(\ram[163][5] ) );
  DFFNX1 \ram_reg[163][4]  ( .D(n2768), .CLK(clk), .Q(\ram[163][4] ) );
  DFFNX1 \ram_reg[163][3]  ( .D(n2767), .CLK(clk), .Q(\ram[163][3] ) );
  DFFNX1 \ram_reg[163][2]  ( .D(n2766), .CLK(clk), .Q(\ram[163][2] ) );
  DFFNX1 \ram_reg[163][1]  ( .D(n2765), .CLK(clk), .Q(\ram[163][1] ) );
  DFFNX1 \ram_reg[163][0]  ( .D(n2764), .CLK(clk), .Q(\ram[163][0] ) );
  DFFNX1 \ram_reg[164][7]  ( .D(n2763), .CLK(clk), .Q(\ram[164][7] ) );
  DFFNX1 \ram_reg[164][6]  ( .D(n2762), .CLK(clk), .Q(\ram[164][6] ) );
  DFFNX1 \ram_reg[164][5]  ( .D(n2761), .CLK(clk), .Q(\ram[164][5] ) );
  DFFNX1 \ram_reg[164][4]  ( .D(n2760), .CLK(clk), .Q(\ram[164][4] ) );
  DFFNX1 \ram_reg[164][3]  ( .D(n2759), .CLK(clk), .Q(\ram[164][3] ) );
  DFFNX1 \ram_reg[164][2]  ( .D(n2758), .CLK(clk), .Q(\ram[164][2] ) );
  DFFNX1 \ram_reg[164][1]  ( .D(n2757), .CLK(clk), .Q(\ram[164][1] ) );
  DFFNX1 \ram_reg[164][0]  ( .D(n2756), .CLK(clk), .Q(\ram[164][0] ) );
  DFFNX1 \ram_reg[165][7]  ( .D(n2755), .CLK(clk), .Q(\ram[165][7] ) );
  DFFNX1 \ram_reg[165][6]  ( .D(n2754), .CLK(clk), .Q(\ram[165][6] ) );
  DFFNX1 \ram_reg[165][5]  ( .D(n2753), .CLK(clk), .Q(\ram[165][5] ) );
  DFFNX1 \ram_reg[165][4]  ( .D(n2752), .CLK(clk), .Q(\ram[165][4] ) );
  DFFNX1 \ram_reg[165][3]  ( .D(n2751), .CLK(clk), .Q(\ram[165][3] ) );
  DFFNX1 \ram_reg[165][2]  ( .D(n2750), .CLK(clk), .Q(\ram[165][2] ) );
  DFFNX1 \ram_reg[165][1]  ( .D(n2749), .CLK(clk), .Q(\ram[165][1] ) );
  DFFNX1 \ram_reg[165][0]  ( .D(n2748), .CLK(clk), .Q(\ram[165][0] ) );
  DFFNX1 \ram_reg[166][7]  ( .D(n2747), .CLK(clk), .Q(\ram[166][7] ) );
  DFFNX1 \ram_reg[166][6]  ( .D(n2746), .CLK(clk), .Q(\ram[166][6] ) );
  DFFNX1 \ram_reg[166][5]  ( .D(n2745), .CLK(clk), .Q(\ram[166][5] ) );
  DFFNX1 \ram_reg[166][4]  ( .D(n2744), .CLK(clk), .Q(\ram[166][4] ) );
  DFFNX1 \ram_reg[166][3]  ( .D(n2743), .CLK(clk), .Q(\ram[166][3] ) );
  DFFNX1 \ram_reg[166][2]  ( .D(n2742), .CLK(clk), .Q(\ram[166][2] ) );
  DFFNX1 \ram_reg[166][1]  ( .D(n2741), .CLK(clk), .Q(\ram[166][1] ) );
  DFFNX1 \ram_reg[166][0]  ( .D(n2740), .CLK(clk), .Q(\ram[166][0] ) );
  DFFNX1 \ram_reg[167][7]  ( .D(n2739), .CLK(clk), .Q(\ram[167][7] ) );
  DFFNX1 \ram_reg[167][6]  ( .D(n2738), .CLK(clk), .Q(\ram[167][6] ) );
  DFFNX1 \ram_reg[167][5]  ( .D(n2737), .CLK(clk), .Q(\ram[167][5] ) );
  DFFNX1 \ram_reg[167][4]  ( .D(n2736), .CLK(clk), .Q(\ram[167][4] ) );
  DFFNX1 \ram_reg[167][3]  ( .D(n2735), .CLK(clk), .Q(\ram[167][3] ) );
  DFFNX1 \ram_reg[167][2]  ( .D(n2734), .CLK(clk), .Q(\ram[167][2] ) );
  DFFNX1 \ram_reg[167][1]  ( .D(n2733), .CLK(clk), .Q(\ram[167][1] ) );
  DFFNX1 \ram_reg[167][0]  ( .D(n2732), .CLK(clk), .Q(\ram[167][0] ) );
  DFFNX1 \ram_reg[168][7]  ( .D(n2731), .CLK(clk), .Q(\ram[168][7] ) );
  DFFNX1 \ram_reg[168][6]  ( .D(n2730), .CLK(clk), .Q(\ram[168][6] ) );
  DFFNX1 \ram_reg[168][5]  ( .D(n2729), .CLK(clk), .Q(\ram[168][5] ) );
  DFFNX1 \ram_reg[168][4]  ( .D(n2728), .CLK(clk), .Q(\ram[168][4] ) );
  DFFNX1 \ram_reg[168][3]  ( .D(n2727), .CLK(clk), .Q(\ram[168][3] ) );
  DFFNX1 \ram_reg[168][2]  ( .D(n2726), .CLK(clk), .Q(\ram[168][2] ) );
  DFFNX1 \ram_reg[168][1]  ( .D(n2725), .CLK(clk), .Q(\ram[168][1] ) );
  DFFNX1 \ram_reg[168][0]  ( .D(n2724), .CLK(clk), .Q(\ram[168][0] ) );
  DFFNX1 \ram_reg[169][7]  ( .D(n2723), .CLK(clk), .Q(\ram[169][7] ) );
  DFFNX1 \ram_reg[169][6]  ( .D(n2722), .CLK(clk), .Q(\ram[169][6] ) );
  DFFNX1 \ram_reg[169][5]  ( .D(n2721), .CLK(clk), .Q(\ram[169][5] ) );
  DFFNX1 \ram_reg[169][4]  ( .D(n2720), .CLK(clk), .Q(\ram[169][4] ) );
  DFFNX1 \ram_reg[169][3]  ( .D(n2719), .CLK(clk), .Q(\ram[169][3] ) );
  DFFNX1 \ram_reg[169][2]  ( .D(n2718), .CLK(clk), .Q(\ram[169][2] ) );
  DFFNX1 \ram_reg[169][1]  ( .D(n2717), .CLK(clk), .Q(\ram[169][1] ) );
  DFFNX1 \ram_reg[169][0]  ( .D(n2716), .CLK(clk), .Q(\ram[169][0] ) );
  DFFNX1 \ram_reg[170][7]  ( .D(n2715), .CLK(clk), .Q(\ram[170][7] ) );
  DFFNX1 \ram_reg[170][6]  ( .D(n2714), .CLK(clk), .Q(\ram[170][6] ) );
  DFFNX1 \ram_reg[170][5]  ( .D(n2713), .CLK(clk), .Q(\ram[170][5] ) );
  DFFNX1 \ram_reg[170][4]  ( .D(n2712), .CLK(clk), .Q(\ram[170][4] ) );
  DFFNX1 \ram_reg[170][3]  ( .D(n2711), .CLK(clk), .Q(\ram[170][3] ) );
  DFFNX1 \ram_reg[170][2]  ( .D(n2710), .CLK(clk), .Q(\ram[170][2] ) );
  DFFNX1 \ram_reg[170][1]  ( .D(n2709), .CLK(clk), .Q(\ram[170][1] ) );
  DFFNX1 \ram_reg[170][0]  ( .D(n2708), .CLK(clk), .Q(\ram[170][0] ) );
  DFFNX1 \ram_reg[171][7]  ( .D(n2707), .CLK(clk), .Q(\ram[171][7] ) );
  DFFNX1 \ram_reg[171][6]  ( .D(n2706), .CLK(clk), .Q(\ram[171][6] ) );
  DFFNX1 \ram_reg[171][5]  ( .D(n2705), .CLK(clk), .Q(\ram[171][5] ) );
  DFFNX1 \ram_reg[171][4]  ( .D(n2704), .CLK(clk), .Q(\ram[171][4] ) );
  DFFNX1 \ram_reg[171][3]  ( .D(n2703), .CLK(clk), .Q(\ram[171][3] ) );
  DFFNX1 \ram_reg[171][2]  ( .D(n2702), .CLK(clk), .Q(\ram[171][2] ) );
  DFFNX1 \ram_reg[171][1]  ( .D(n2701), .CLK(clk), .Q(\ram[171][1] ) );
  DFFNX1 \ram_reg[171][0]  ( .D(n2700), .CLK(clk), .Q(\ram[171][0] ) );
  DFFNX1 \ram_reg[172][7]  ( .D(n2699), .CLK(clk), .Q(\ram[172][7] ) );
  DFFNX1 \ram_reg[172][6]  ( .D(n2698), .CLK(clk), .Q(\ram[172][6] ) );
  DFFNX1 \ram_reg[172][5]  ( .D(n2697), .CLK(clk), .Q(\ram[172][5] ) );
  DFFNX1 \ram_reg[172][4]  ( .D(n2696), .CLK(clk), .Q(\ram[172][4] ) );
  DFFNX1 \ram_reg[172][3]  ( .D(n2695), .CLK(clk), .Q(\ram[172][3] ) );
  DFFNX1 \ram_reg[172][2]  ( .D(n2694), .CLK(clk), .Q(\ram[172][2] ) );
  DFFNX1 \ram_reg[172][1]  ( .D(n2693), .CLK(clk), .Q(\ram[172][1] ) );
  DFFNX1 \ram_reg[172][0]  ( .D(n2692), .CLK(clk), .Q(\ram[172][0] ) );
  DFFNX1 \ram_reg[173][7]  ( .D(n2691), .CLK(clk), .Q(\ram[173][7] ) );
  DFFNX1 \ram_reg[173][6]  ( .D(n2690), .CLK(clk), .Q(\ram[173][6] ) );
  DFFNX1 \ram_reg[173][5]  ( .D(n2689), .CLK(clk), .Q(\ram[173][5] ) );
  DFFNX1 \ram_reg[173][4]  ( .D(n2688), .CLK(clk), .Q(\ram[173][4] ) );
  DFFNX1 \ram_reg[173][3]  ( .D(n2687), .CLK(clk), .Q(\ram[173][3] ) );
  DFFNX1 \ram_reg[173][2]  ( .D(n2686), .CLK(clk), .Q(\ram[173][2] ) );
  DFFNX1 \ram_reg[173][1]  ( .D(n2685), .CLK(clk), .Q(\ram[173][1] ) );
  DFFNX1 \ram_reg[173][0]  ( .D(n2684), .CLK(clk), .Q(\ram[173][0] ) );
  DFFNX1 \ram_reg[174][7]  ( .D(n2683), .CLK(clk), .Q(\ram[174][7] ) );
  DFFNX1 \ram_reg[174][6]  ( .D(n2682), .CLK(clk), .Q(\ram[174][6] ) );
  DFFNX1 \ram_reg[174][5]  ( .D(n2681), .CLK(clk), .Q(\ram[174][5] ) );
  DFFNX1 \ram_reg[174][4]  ( .D(n2680), .CLK(clk), .Q(\ram[174][4] ) );
  DFFNX1 \ram_reg[174][3]  ( .D(n2679), .CLK(clk), .Q(\ram[174][3] ) );
  DFFNX1 \ram_reg[174][2]  ( .D(n2678), .CLK(clk), .Q(\ram[174][2] ) );
  DFFNX1 \ram_reg[174][1]  ( .D(n2677), .CLK(clk), .Q(\ram[174][1] ) );
  DFFNX1 \ram_reg[174][0]  ( .D(n2676), .CLK(clk), .Q(\ram[174][0] ) );
  DFFNX1 \ram_reg[175][7]  ( .D(n2675), .CLK(clk), .Q(\ram[175][7] ) );
  DFFNX1 \ram_reg[175][6]  ( .D(n2674), .CLK(clk), .Q(\ram[175][6] ) );
  DFFNX1 \ram_reg[175][5]  ( .D(n2673), .CLK(clk), .Q(\ram[175][5] ) );
  DFFNX1 \ram_reg[175][4]  ( .D(n2672), .CLK(clk), .Q(\ram[175][4] ) );
  DFFNX1 \ram_reg[175][3]  ( .D(n2671), .CLK(clk), .Q(\ram[175][3] ) );
  DFFNX1 \ram_reg[175][2]  ( .D(n2670), .CLK(clk), .Q(\ram[175][2] ) );
  DFFNX1 \ram_reg[175][1]  ( .D(n2669), .CLK(clk), .Q(\ram[175][1] ) );
  DFFNX1 \ram_reg[175][0]  ( .D(n2668), .CLK(clk), .Q(\ram[175][0] ) );
  DFFNX1 \ram_reg[176][7]  ( .D(n2667), .CLK(clk), .Q(\ram[176][7] ) );
  DFFNX1 \ram_reg[176][6]  ( .D(n2666), .CLK(clk), .Q(\ram[176][6] ) );
  DFFNX1 \ram_reg[176][5]  ( .D(n2665), .CLK(clk), .Q(\ram[176][5] ) );
  DFFNX1 \ram_reg[176][4]  ( .D(n2664), .CLK(clk), .Q(\ram[176][4] ) );
  DFFNX1 \ram_reg[176][3]  ( .D(n2663), .CLK(clk), .Q(\ram[176][3] ) );
  DFFNX1 \ram_reg[176][2]  ( .D(n2662), .CLK(clk), .Q(\ram[176][2] ) );
  DFFNX1 \ram_reg[176][1]  ( .D(n2661), .CLK(clk), .Q(\ram[176][1] ) );
  DFFNX1 \ram_reg[176][0]  ( .D(n2660), .CLK(clk), .Q(\ram[176][0] ) );
  DFFNX1 \ram_reg[177][7]  ( .D(n2659), .CLK(clk), .Q(\ram[177][7] ) );
  DFFNX1 \ram_reg[177][6]  ( .D(n2658), .CLK(clk), .Q(\ram[177][6] ) );
  DFFNX1 \ram_reg[177][5]  ( .D(n2657), .CLK(clk), .Q(\ram[177][5] ) );
  DFFNX1 \ram_reg[177][4]  ( .D(n2656), .CLK(clk), .Q(\ram[177][4] ) );
  DFFNX1 \ram_reg[177][3]  ( .D(n2655), .CLK(clk), .Q(\ram[177][3] ) );
  DFFNX1 \ram_reg[177][2]  ( .D(n2654), .CLK(clk), .Q(\ram[177][2] ) );
  DFFNX1 \ram_reg[177][1]  ( .D(n2653), .CLK(clk), .Q(\ram[177][1] ) );
  DFFNX1 \ram_reg[177][0]  ( .D(n2652), .CLK(clk), .Q(\ram[177][0] ) );
  DFFNX1 \ram_reg[178][7]  ( .D(n2651), .CLK(clk), .Q(\ram[178][7] ) );
  DFFNX1 \ram_reg[178][6]  ( .D(n2650), .CLK(clk), .Q(\ram[178][6] ) );
  DFFNX1 \ram_reg[178][5]  ( .D(n2649), .CLK(clk), .Q(\ram[178][5] ) );
  DFFNX1 \ram_reg[178][4]  ( .D(n2648), .CLK(clk), .Q(\ram[178][4] ) );
  DFFNX1 \ram_reg[178][3]  ( .D(n2647), .CLK(clk), .Q(\ram[178][3] ) );
  DFFNX1 \ram_reg[178][2]  ( .D(n2646), .CLK(clk), .Q(\ram[178][2] ) );
  DFFNX1 \ram_reg[178][1]  ( .D(n2645), .CLK(clk), .Q(\ram[178][1] ) );
  DFFNX1 \ram_reg[178][0]  ( .D(n2644), .CLK(clk), .Q(\ram[178][0] ) );
  DFFNX1 \ram_reg[179][7]  ( .D(n2643), .CLK(clk), .Q(\ram[179][7] ) );
  DFFNX1 \ram_reg[179][6]  ( .D(n2642), .CLK(clk), .Q(\ram[179][6] ) );
  DFFNX1 \ram_reg[179][5]  ( .D(n2641), .CLK(clk), .Q(\ram[179][5] ) );
  DFFNX1 \ram_reg[179][4]  ( .D(n2640), .CLK(clk), .Q(\ram[179][4] ) );
  DFFNX1 \ram_reg[179][3]  ( .D(n2639), .CLK(clk), .Q(\ram[179][3] ) );
  DFFNX1 \ram_reg[179][2]  ( .D(n2638), .CLK(clk), .Q(\ram[179][2] ) );
  DFFNX1 \ram_reg[179][1]  ( .D(n2637), .CLK(clk), .Q(\ram[179][1] ) );
  DFFNX1 \ram_reg[179][0]  ( .D(n2636), .CLK(clk), .Q(\ram[179][0] ) );
  DFFNX1 \ram_reg[180][7]  ( .D(n2635), .CLK(clk), .Q(\ram[180][7] ) );
  DFFNX1 \ram_reg[180][6]  ( .D(n2634), .CLK(clk), .Q(\ram[180][6] ) );
  DFFNX1 \ram_reg[180][5]  ( .D(n2633), .CLK(clk), .Q(\ram[180][5] ) );
  DFFNX1 \ram_reg[180][4]  ( .D(n2632), .CLK(clk), .Q(\ram[180][4] ) );
  DFFNX1 \ram_reg[180][3]  ( .D(n2631), .CLK(clk), .Q(\ram[180][3] ) );
  DFFNX1 \ram_reg[180][2]  ( .D(n2630), .CLK(clk), .Q(\ram[180][2] ) );
  DFFNX1 \ram_reg[180][1]  ( .D(n2629), .CLK(clk), .Q(\ram[180][1] ) );
  DFFNX1 \ram_reg[180][0]  ( .D(n2628), .CLK(clk), .Q(\ram[180][0] ) );
  DFFNX1 \ram_reg[181][7]  ( .D(n2627), .CLK(clk), .Q(\ram[181][7] ) );
  DFFNX1 \ram_reg[181][6]  ( .D(n2626), .CLK(clk), .Q(\ram[181][6] ) );
  DFFNX1 \ram_reg[181][5]  ( .D(n2625), .CLK(clk), .Q(\ram[181][5] ) );
  DFFNX1 \ram_reg[181][4]  ( .D(n2624), .CLK(clk), .Q(\ram[181][4] ) );
  DFFNX1 \ram_reg[181][3]  ( .D(n2623), .CLK(clk), .Q(\ram[181][3] ) );
  DFFNX1 \ram_reg[181][2]  ( .D(n2622), .CLK(clk), .Q(\ram[181][2] ) );
  DFFNX1 \ram_reg[181][1]  ( .D(n2621), .CLK(clk), .Q(\ram[181][1] ) );
  DFFNX1 \ram_reg[181][0]  ( .D(n2620), .CLK(clk), .Q(\ram[181][0] ) );
  DFFNX1 \ram_reg[182][7]  ( .D(n2619), .CLK(clk), .Q(\ram[182][7] ) );
  DFFNX1 \ram_reg[182][6]  ( .D(n2618), .CLK(clk), .Q(\ram[182][6] ) );
  DFFNX1 \ram_reg[182][5]  ( .D(n2617), .CLK(clk), .Q(\ram[182][5] ) );
  DFFNX1 \ram_reg[182][4]  ( .D(n2616), .CLK(clk), .Q(\ram[182][4] ) );
  DFFNX1 \ram_reg[182][3]  ( .D(n2615), .CLK(clk), .Q(\ram[182][3] ) );
  DFFNX1 \ram_reg[182][2]  ( .D(n2614), .CLK(clk), .Q(\ram[182][2] ) );
  DFFNX1 \ram_reg[182][1]  ( .D(n2613), .CLK(clk), .Q(\ram[182][1] ) );
  DFFNX1 \ram_reg[182][0]  ( .D(n2612), .CLK(clk), .Q(\ram[182][0] ) );
  DFFNX1 \ram_reg[183][7]  ( .D(n2611), .CLK(clk), .Q(\ram[183][7] ) );
  DFFNX1 \ram_reg[183][6]  ( .D(n2610), .CLK(clk), .Q(\ram[183][6] ) );
  DFFNX1 \ram_reg[183][5]  ( .D(n2609), .CLK(clk), .Q(\ram[183][5] ) );
  DFFNX1 \ram_reg[183][4]  ( .D(n2608), .CLK(clk), .Q(\ram[183][4] ) );
  DFFNX1 \ram_reg[183][3]  ( .D(n2607), .CLK(clk), .Q(\ram[183][3] ) );
  DFFNX1 \ram_reg[183][2]  ( .D(n2606), .CLK(clk), .Q(\ram[183][2] ) );
  DFFNX1 \ram_reg[183][1]  ( .D(n2605), .CLK(clk), .Q(\ram[183][1] ) );
  DFFNX1 \ram_reg[183][0]  ( .D(n2604), .CLK(clk), .Q(\ram[183][0] ) );
  DFFNX1 \ram_reg[184][7]  ( .D(n2603), .CLK(clk), .Q(\ram[184][7] ) );
  DFFNX1 \ram_reg[184][6]  ( .D(n2602), .CLK(clk), .Q(\ram[184][6] ) );
  DFFNX1 \ram_reg[184][5]  ( .D(n2601), .CLK(clk), .Q(\ram[184][5] ) );
  DFFNX1 \ram_reg[184][4]  ( .D(n2600), .CLK(clk), .Q(\ram[184][4] ) );
  DFFNX1 \ram_reg[184][3]  ( .D(n2599), .CLK(clk), .Q(\ram[184][3] ) );
  DFFNX1 \ram_reg[184][2]  ( .D(n2598), .CLK(clk), .Q(\ram[184][2] ) );
  DFFNX1 \ram_reg[184][1]  ( .D(n2597), .CLK(clk), .Q(\ram[184][1] ) );
  DFFNX1 \ram_reg[184][0]  ( .D(n2596), .CLK(clk), .Q(\ram[184][0] ) );
  DFFNX1 \ram_reg[185][7]  ( .D(n2595), .CLK(clk), .Q(\ram[185][7] ) );
  DFFNX1 \ram_reg[185][6]  ( .D(n2594), .CLK(clk), .Q(\ram[185][6] ) );
  DFFNX1 \ram_reg[185][5]  ( .D(n2593), .CLK(clk), .Q(\ram[185][5] ) );
  DFFNX1 \ram_reg[185][4]  ( .D(n2592), .CLK(clk), .Q(\ram[185][4] ) );
  DFFNX1 \ram_reg[185][3]  ( .D(n2591), .CLK(clk), .Q(\ram[185][3] ) );
  DFFNX1 \ram_reg[185][2]  ( .D(n2590), .CLK(clk), .Q(\ram[185][2] ) );
  DFFNX1 \ram_reg[185][1]  ( .D(n2589), .CLK(clk), .Q(\ram[185][1] ) );
  DFFNX1 \ram_reg[185][0]  ( .D(n2588), .CLK(clk), .Q(\ram[185][0] ) );
  DFFNX1 \ram_reg[186][7]  ( .D(n2587), .CLK(clk), .Q(\ram[186][7] ) );
  DFFNX1 \ram_reg[186][6]  ( .D(n2586), .CLK(clk), .Q(\ram[186][6] ) );
  DFFNX1 \ram_reg[186][5]  ( .D(n2585), .CLK(clk), .Q(\ram[186][5] ) );
  DFFNX1 \ram_reg[186][4]  ( .D(n2584), .CLK(clk), .Q(\ram[186][4] ) );
  DFFNX1 \ram_reg[186][3]  ( .D(n2583), .CLK(clk), .Q(\ram[186][3] ) );
  DFFNX1 \ram_reg[186][2]  ( .D(n2582), .CLK(clk), .Q(\ram[186][2] ) );
  DFFNX1 \ram_reg[186][1]  ( .D(n2581), .CLK(clk), .Q(\ram[186][1] ) );
  DFFNX1 \ram_reg[186][0]  ( .D(n2580), .CLK(clk), .Q(\ram[186][0] ) );
  DFFNX1 \ram_reg[187][7]  ( .D(n2579), .CLK(clk), .Q(\ram[187][7] ) );
  DFFNX1 \ram_reg[187][6]  ( .D(n2578), .CLK(clk), .Q(\ram[187][6] ) );
  DFFNX1 \ram_reg[187][5]  ( .D(n2577), .CLK(clk), .Q(\ram[187][5] ) );
  DFFNX1 \ram_reg[187][4]  ( .D(n2576), .CLK(clk), .Q(\ram[187][4] ) );
  DFFNX1 \ram_reg[187][3]  ( .D(n2575), .CLK(clk), .Q(\ram[187][3] ) );
  DFFNX1 \ram_reg[187][2]  ( .D(n2574), .CLK(clk), .Q(\ram[187][2] ) );
  DFFNX1 \ram_reg[187][1]  ( .D(n2573), .CLK(clk), .Q(\ram[187][1] ) );
  DFFNX1 \ram_reg[187][0]  ( .D(n2572), .CLK(clk), .Q(\ram[187][0] ) );
  DFFNX1 \ram_reg[188][7]  ( .D(n2571), .CLK(clk), .Q(\ram[188][7] ) );
  DFFNX1 \ram_reg[188][6]  ( .D(n2570), .CLK(clk), .Q(\ram[188][6] ) );
  DFFNX1 \ram_reg[188][5]  ( .D(n2569), .CLK(clk), .Q(\ram[188][5] ) );
  DFFNX1 \ram_reg[188][4]  ( .D(n2568), .CLK(clk), .Q(\ram[188][4] ) );
  DFFNX1 \ram_reg[188][3]  ( .D(n2567), .CLK(clk), .Q(\ram[188][3] ) );
  DFFNX1 \ram_reg[188][2]  ( .D(n2566), .CLK(clk), .Q(\ram[188][2] ) );
  DFFNX1 \ram_reg[188][1]  ( .D(n2565), .CLK(clk), .Q(\ram[188][1] ) );
  DFFNX1 \ram_reg[188][0]  ( .D(n2564), .CLK(clk), .Q(\ram[188][0] ) );
  DFFNX1 \ram_reg[189][7]  ( .D(n2563), .CLK(clk), .Q(\ram[189][7] ) );
  DFFNX1 \ram_reg[189][6]  ( .D(n2562), .CLK(clk), .Q(\ram[189][6] ) );
  DFFNX1 \ram_reg[189][5]  ( .D(n2561), .CLK(clk), .Q(\ram[189][5] ) );
  DFFNX1 \ram_reg[189][4]  ( .D(n2560), .CLK(clk), .Q(\ram[189][4] ) );
  DFFNX1 \ram_reg[189][3]  ( .D(n2559), .CLK(clk), .Q(\ram[189][3] ) );
  DFFNX1 \ram_reg[189][2]  ( .D(n2558), .CLK(clk), .Q(\ram[189][2] ) );
  DFFNX1 \ram_reg[189][1]  ( .D(n2557), .CLK(clk), .Q(\ram[189][1] ) );
  DFFNX1 \ram_reg[189][0]  ( .D(n2556), .CLK(clk), .Q(\ram[189][0] ) );
  DFFNX1 \ram_reg[190][7]  ( .D(n2555), .CLK(clk), .Q(\ram[190][7] ) );
  DFFNX1 \ram_reg[190][6]  ( .D(n2554), .CLK(clk), .Q(\ram[190][6] ) );
  DFFNX1 \ram_reg[190][5]  ( .D(n2553), .CLK(clk), .Q(\ram[190][5] ) );
  DFFNX1 \ram_reg[190][4]  ( .D(n2552), .CLK(clk), .Q(\ram[190][4] ) );
  DFFNX1 \ram_reg[190][3]  ( .D(n2551), .CLK(clk), .Q(\ram[190][3] ) );
  DFFNX1 \ram_reg[190][2]  ( .D(n2550), .CLK(clk), .Q(\ram[190][2] ) );
  DFFNX1 \ram_reg[190][1]  ( .D(n2549), .CLK(clk), .Q(\ram[190][1] ) );
  DFFNX1 \ram_reg[190][0]  ( .D(n2548), .CLK(clk), .Q(\ram[190][0] ) );
  DFFNX1 \ram_reg[191][7]  ( .D(n2547), .CLK(clk), .Q(\ram[191][7] ) );
  DFFNX1 \ram_reg[191][6]  ( .D(n2546), .CLK(clk), .Q(\ram[191][6] ) );
  DFFNX1 \ram_reg[191][5]  ( .D(n2545), .CLK(clk), .Q(\ram[191][5] ) );
  DFFNX1 \ram_reg[191][4]  ( .D(n2544), .CLK(clk), .Q(\ram[191][4] ) );
  DFFNX1 \ram_reg[191][3]  ( .D(n2543), .CLK(clk), .Q(\ram[191][3] ) );
  DFFNX1 \ram_reg[191][2]  ( .D(n2542), .CLK(clk), .Q(\ram[191][2] ) );
  DFFNX1 \ram_reg[191][1]  ( .D(n2541), .CLK(clk), .Q(\ram[191][1] ) );
  DFFNX1 \ram_reg[191][0]  ( .D(n2540), .CLK(clk), .Q(\ram[191][0] ) );
  DFFNX1 \ram_reg[192][7]  ( .D(n2539), .CLK(clk), .Q(\ram[192][7] ) );
  DFFNX1 \ram_reg[192][6]  ( .D(n2538), .CLK(clk), .Q(\ram[192][6] ) );
  DFFNX1 \ram_reg[192][5]  ( .D(n2537), .CLK(clk), .Q(\ram[192][5] ) );
  DFFNX1 \ram_reg[192][4]  ( .D(n2536), .CLK(clk), .Q(\ram[192][4] ) );
  DFFNX1 \ram_reg[192][3]  ( .D(n2535), .CLK(clk), .Q(\ram[192][3] ) );
  DFFNX1 \ram_reg[192][2]  ( .D(n2534), .CLK(clk), .Q(\ram[192][2] ) );
  DFFNX1 \ram_reg[192][1]  ( .D(n2533), .CLK(clk), .Q(\ram[192][1] ) );
  DFFNX1 \ram_reg[192][0]  ( .D(n2532), .CLK(clk), .Q(\ram[192][0] ) );
  DFFNX1 \ram_reg[193][7]  ( .D(n2531), .CLK(clk), .Q(\ram[193][7] ) );
  DFFNX1 \ram_reg[193][6]  ( .D(n2530), .CLK(clk), .Q(\ram[193][6] ) );
  DFFNX1 \ram_reg[193][5]  ( .D(n2529), .CLK(clk), .Q(\ram[193][5] ) );
  DFFNX1 \ram_reg[193][4]  ( .D(n2528), .CLK(clk), .Q(\ram[193][4] ) );
  DFFNX1 \ram_reg[193][3]  ( .D(n2527), .CLK(clk), .Q(\ram[193][3] ) );
  DFFNX1 \ram_reg[193][2]  ( .D(n2526), .CLK(clk), .Q(\ram[193][2] ) );
  DFFNX1 \ram_reg[193][1]  ( .D(n2525), .CLK(clk), .Q(\ram[193][1] ) );
  DFFNX1 \ram_reg[193][0]  ( .D(n2524), .CLK(clk), .Q(\ram[193][0] ) );
  DFFNX1 \ram_reg[194][7]  ( .D(n2523), .CLK(clk), .Q(\ram[194][7] ) );
  DFFNX1 \ram_reg[194][6]  ( .D(n2522), .CLK(clk), .Q(\ram[194][6] ) );
  DFFNX1 \ram_reg[194][5]  ( .D(n2521), .CLK(clk), .Q(\ram[194][5] ) );
  DFFNX1 \ram_reg[194][4]  ( .D(n2520), .CLK(clk), .Q(\ram[194][4] ) );
  DFFNX1 \ram_reg[194][3]  ( .D(n2519), .CLK(clk), .Q(\ram[194][3] ) );
  DFFNX1 \ram_reg[194][2]  ( .D(n2518), .CLK(clk), .Q(\ram[194][2] ) );
  DFFNX1 \ram_reg[194][1]  ( .D(n2517), .CLK(clk), .Q(\ram[194][1] ) );
  DFFNX1 \ram_reg[194][0]  ( .D(n2516), .CLK(clk), .Q(\ram[194][0] ) );
  DFFNX1 \ram_reg[195][7]  ( .D(n2515), .CLK(clk), .Q(\ram[195][7] ) );
  DFFNX1 \ram_reg[195][6]  ( .D(n2514), .CLK(clk), .Q(\ram[195][6] ) );
  DFFNX1 \ram_reg[195][5]  ( .D(n2513), .CLK(clk), .Q(\ram[195][5] ) );
  DFFNX1 \ram_reg[195][4]  ( .D(n2512), .CLK(clk), .Q(\ram[195][4] ) );
  DFFNX1 \ram_reg[195][3]  ( .D(n2511), .CLK(clk), .Q(\ram[195][3] ) );
  DFFNX1 \ram_reg[195][2]  ( .D(n2510), .CLK(clk), .Q(\ram[195][2] ) );
  DFFNX1 \ram_reg[195][1]  ( .D(n2509), .CLK(clk), .Q(\ram[195][1] ) );
  DFFNX1 \ram_reg[195][0]  ( .D(n2508), .CLK(clk), .Q(\ram[195][0] ) );
  DFFNX1 \ram_reg[196][7]  ( .D(n2507), .CLK(clk), .Q(\ram[196][7] ) );
  DFFNX1 \ram_reg[196][6]  ( .D(n2506), .CLK(clk), .Q(\ram[196][6] ) );
  DFFNX1 \ram_reg[196][5]  ( .D(n2505), .CLK(clk), .Q(\ram[196][5] ) );
  DFFNX1 \ram_reg[196][4]  ( .D(n2504), .CLK(clk), .Q(\ram[196][4] ) );
  DFFNX1 \ram_reg[196][3]  ( .D(n2503), .CLK(clk), .Q(\ram[196][3] ) );
  DFFNX1 \ram_reg[196][2]  ( .D(n2502), .CLK(clk), .Q(\ram[196][2] ) );
  DFFNX1 \ram_reg[196][1]  ( .D(n2501), .CLK(clk), .Q(\ram[196][1] ) );
  DFFNX1 \ram_reg[196][0]  ( .D(n2500), .CLK(clk), .Q(\ram[196][0] ) );
  DFFNX1 \ram_reg[197][7]  ( .D(n2499), .CLK(clk), .Q(\ram[197][7] ) );
  DFFNX1 \ram_reg[197][6]  ( .D(n2498), .CLK(clk), .Q(\ram[197][6] ) );
  DFFNX1 \ram_reg[197][5]  ( .D(n2497), .CLK(clk), .Q(\ram[197][5] ) );
  DFFNX1 \ram_reg[197][4]  ( .D(n2496), .CLK(clk), .Q(\ram[197][4] ) );
  DFFNX1 \ram_reg[197][3]  ( .D(n2495), .CLK(clk), .Q(\ram[197][3] ) );
  DFFNX1 \ram_reg[197][2]  ( .D(n2494), .CLK(clk), .Q(\ram[197][2] ) );
  DFFNX1 \ram_reg[197][1]  ( .D(n2493), .CLK(clk), .Q(\ram[197][1] ) );
  DFFNX1 \ram_reg[197][0]  ( .D(n2492), .CLK(clk), .Q(\ram[197][0] ) );
  DFFNX1 \ram_reg[198][7]  ( .D(n2491), .CLK(clk), .Q(\ram[198][7] ) );
  DFFNX1 \ram_reg[198][6]  ( .D(n2490), .CLK(clk), .Q(\ram[198][6] ) );
  DFFNX1 \ram_reg[198][5]  ( .D(n2489), .CLK(clk), .Q(\ram[198][5] ) );
  DFFNX1 \ram_reg[198][4]  ( .D(n2488), .CLK(clk), .Q(\ram[198][4] ) );
  DFFNX1 \ram_reg[198][3]  ( .D(n2487), .CLK(clk), .Q(\ram[198][3] ) );
  DFFNX1 \ram_reg[198][2]  ( .D(n2486), .CLK(clk), .Q(\ram[198][2] ) );
  DFFNX1 \ram_reg[198][1]  ( .D(n2485), .CLK(clk), .Q(\ram[198][1] ) );
  DFFNX1 \ram_reg[198][0]  ( .D(n2484), .CLK(clk), .Q(\ram[198][0] ) );
  DFFNX1 \ram_reg[199][7]  ( .D(n2483), .CLK(clk), .Q(\ram[199][7] ) );
  DFFNX1 \ram_reg[199][6]  ( .D(n2482), .CLK(clk), .Q(\ram[199][6] ) );
  DFFNX1 \ram_reg[199][5]  ( .D(n2481), .CLK(clk), .Q(\ram[199][5] ) );
  DFFNX1 \ram_reg[199][4]  ( .D(n2480), .CLK(clk), .Q(\ram[199][4] ) );
  DFFNX1 \ram_reg[199][3]  ( .D(n2479), .CLK(clk), .Q(\ram[199][3] ) );
  DFFNX1 \ram_reg[199][2]  ( .D(n2478), .CLK(clk), .Q(\ram[199][2] ) );
  DFFNX1 \ram_reg[199][1]  ( .D(n2477), .CLK(clk), .Q(\ram[199][1] ) );
  DFFNX1 \ram_reg[199][0]  ( .D(n2476), .CLK(clk), .Q(\ram[199][0] ) );
  DFFNX1 \ram_reg[200][7]  ( .D(n2475), .CLK(clk), .Q(\ram[200][7] ) );
  DFFNX1 \ram_reg[200][6]  ( .D(n2474), .CLK(clk), .Q(\ram[200][6] ) );
  DFFNX1 \ram_reg[200][5]  ( .D(n2473), .CLK(clk), .Q(\ram[200][5] ) );
  DFFNX1 \ram_reg[200][4]  ( .D(n2472), .CLK(clk), .Q(\ram[200][4] ) );
  DFFNX1 \ram_reg[200][3]  ( .D(n2471), .CLK(clk), .Q(\ram[200][3] ) );
  DFFNX1 \ram_reg[200][2]  ( .D(n2470), .CLK(clk), .Q(\ram[200][2] ) );
  DFFNX1 \ram_reg[200][1]  ( .D(n2469), .CLK(clk), .Q(\ram[200][1] ) );
  DFFNX1 \ram_reg[200][0]  ( .D(n2468), .CLK(clk), .Q(\ram[200][0] ) );
  DFFNX1 \ram_reg[201][7]  ( .D(n2467), .CLK(clk), .Q(\ram[201][7] ) );
  DFFNX1 \ram_reg[201][6]  ( .D(n2466), .CLK(clk), .Q(\ram[201][6] ) );
  DFFNX1 \ram_reg[201][5]  ( .D(n2465), .CLK(clk), .Q(\ram[201][5] ) );
  DFFNX1 \ram_reg[201][4]  ( .D(n2464), .CLK(clk), .Q(\ram[201][4] ) );
  DFFNX1 \ram_reg[201][3]  ( .D(n2463), .CLK(clk), .Q(\ram[201][3] ) );
  DFFNX1 \ram_reg[201][2]  ( .D(n2462), .CLK(clk), .Q(\ram[201][2] ) );
  DFFNX1 \ram_reg[201][1]  ( .D(n2461), .CLK(clk), .Q(\ram[201][1] ) );
  DFFNX1 \ram_reg[201][0]  ( .D(n2460), .CLK(clk), .Q(\ram[201][0] ) );
  DFFNX1 \ram_reg[202][7]  ( .D(n2459), .CLK(clk), .Q(\ram[202][7] ) );
  DFFNX1 \ram_reg[202][6]  ( .D(n2458), .CLK(clk), .Q(\ram[202][6] ) );
  DFFNX1 \ram_reg[202][5]  ( .D(n2457), .CLK(clk), .Q(\ram[202][5] ) );
  DFFNX1 \ram_reg[202][4]  ( .D(n2456), .CLK(clk), .Q(\ram[202][4] ) );
  DFFNX1 \ram_reg[202][3]  ( .D(n2455), .CLK(clk), .Q(\ram[202][3] ) );
  DFFNX1 \ram_reg[202][2]  ( .D(n2454), .CLK(clk), .Q(\ram[202][2] ) );
  DFFNX1 \ram_reg[202][1]  ( .D(n2453), .CLK(clk), .Q(\ram[202][1] ) );
  DFFNX1 \ram_reg[202][0]  ( .D(n2452), .CLK(clk), .Q(\ram[202][0] ) );
  DFFNX1 \ram_reg[203][7]  ( .D(n2451), .CLK(clk), .Q(\ram[203][7] ) );
  DFFNX1 \ram_reg[203][6]  ( .D(n2450), .CLK(clk), .Q(\ram[203][6] ) );
  DFFNX1 \ram_reg[203][5]  ( .D(n2449), .CLK(clk), .Q(\ram[203][5] ) );
  DFFNX1 \ram_reg[203][4]  ( .D(n2448), .CLK(clk), .Q(\ram[203][4] ) );
  DFFNX1 \ram_reg[203][3]  ( .D(n2447), .CLK(clk), .Q(\ram[203][3] ) );
  DFFNX1 \ram_reg[203][2]  ( .D(n2446), .CLK(clk), .Q(\ram[203][2] ) );
  DFFNX1 \ram_reg[203][1]  ( .D(n2445), .CLK(clk), .Q(\ram[203][1] ) );
  DFFNX1 \ram_reg[203][0]  ( .D(n2444), .CLK(clk), .Q(\ram[203][0] ) );
  DFFNX1 \ram_reg[204][7]  ( .D(n2443), .CLK(clk), .Q(\ram[204][7] ) );
  DFFNX1 \ram_reg[204][6]  ( .D(n2442), .CLK(clk), .Q(\ram[204][6] ) );
  DFFNX1 \ram_reg[204][5]  ( .D(n2441), .CLK(clk), .Q(\ram[204][5] ) );
  DFFNX1 \ram_reg[204][4]  ( .D(n2440), .CLK(clk), .Q(\ram[204][4] ) );
  DFFNX1 \ram_reg[204][3]  ( .D(n2439), .CLK(clk), .Q(\ram[204][3] ) );
  DFFNX1 \ram_reg[204][2]  ( .D(n2438), .CLK(clk), .Q(\ram[204][2] ) );
  DFFNX1 \ram_reg[204][1]  ( .D(n2437), .CLK(clk), .Q(\ram[204][1] ) );
  DFFNX1 \ram_reg[204][0]  ( .D(n2436), .CLK(clk), .Q(\ram[204][0] ) );
  DFFNX1 \ram_reg[205][7]  ( .D(n2435), .CLK(clk), .Q(\ram[205][7] ) );
  DFFNX1 \ram_reg[205][6]  ( .D(n2434), .CLK(clk), .Q(\ram[205][6] ) );
  DFFNX1 \ram_reg[205][5]  ( .D(n2433), .CLK(clk), .Q(\ram[205][5] ) );
  DFFNX1 \ram_reg[205][4]  ( .D(n2432), .CLK(clk), .Q(\ram[205][4] ) );
  DFFNX1 \ram_reg[205][3]  ( .D(n2431), .CLK(clk), .Q(\ram[205][3] ) );
  DFFNX1 \ram_reg[205][2]  ( .D(n2430), .CLK(clk), .Q(\ram[205][2] ) );
  DFFNX1 \ram_reg[205][1]  ( .D(n2429), .CLK(clk), .Q(\ram[205][1] ) );
  DFFNX1 \ram_reg[205][0]  ( .D(n2428), .CLK(clk), .Q(\ram[205][0] ) );
  DFFNX1 \ram_reg[206][7]  ( .D(n2427), .CLK(clk), .Q(\ram[206][7] ) );
  DFFNX1 \ram_reg[206][6]  ( .D(n2426), .CLK(clk), .Q(\ram[206][6] ) );
  DFFNX1 \ram_reg[206][5]  ( .D(n2425), .CLK(clk), .Q(\ram[206][5] ) );
  DFFNX1 \ram_reg[206][4]  ( .D(n2424), .CLK(clk), .Q(\ram[206][4] ) );
  DFFNX1 \ram_reg[206][3]  ( .D(n2423), .CLK(clk), .Q(\ram[206][3] ) );
  DFFNX1 \ram_reg[206][2]  ( .D(n2422), .CLK(clk), .Q(\ram[206][2] ) );
  DFFNX1 \ram_reg[206][1]  ( .D(n2421), .CLK(clk), .Q(\ram[206][1] ) );
  DFFNX1 \ram_reg[206][0]  ( .D(n2420), .CLK(clk), .Q(\ram[206][0] ) );
  DFFNX1 \ram_reg[207][7]  ( .D(n2419), .CLK(clk), .Q(\ram[207][7] ) );
  DFFNX1 \ram_reg[207][6]  ( .D(n2418), .CLK(clk), .Q(\ram[207][6] ) );
  DFFNX1 \ram_reg[207][5]  ( .D(n2417), .CLK(clk), .Q(\ram[207][5] ) );
  DFFNX1 \ram_reg[207][4]  ( .D(n2416), .CLK(clk), .Q(\ram[207][4] ) );
  DFFNX1 \ram_reg[207][3]  ( .D(n2415), .CLK(clk), .Q(\ram[207][3] ) );
  DFFNX1 \ram_reg[207][2]  ( .D(n2414), .CLK(clk), .Q(\ram[207][2] ) );
  DFFNX1 \ram_reg[207][1]  ( .D(n2413), .CLK(clk), .Q(\ram[207][1] ) );
  DFFNX1 \ram_reg[207][0]  ( .D(n2412), .CLK(clk), .Q(\ram[207][0] ) );
  DFFNX1 \ram_reg[208][7]  ( .D(n2411), .CLK(clk), .Q(\ram[208][7] ) );
  DFFNX1 \ram_reg[208][6]  ( .D(n2410), .CLK(clk), .Q(\ram[208][6] ) );
  DFFNX1 \ram_reg[208][5]  ( .D(n2409), .CLK(clk), .Q(\ram[208][5] ) );
  DFFNX1 \ram_reg[208][4]  ( .D(n2408), .CLK(clk), .Q(\ram[208][4] ) );
  DFFNX1 \ram_reg[208][3]  ( .D(n2407), .CLK(clk), .Q(\ram[208][3] ) );
  DFFNX1 \ram_reg[208][2]  ( .D(n2406), .CLK(clk), .Q(\ram[208][2] ) );
  DFFNX1 \ram_reg[208][1]  ( .D(n2405), .CLK(clk), .Q(\ram[208][1] ) );
  DFFNX1 \ram_reg[208][0]  ( .D(n2404), .CLK(clk), .Q(\ram[208][0] ) );
  DFFNX1 \ram_reg[209][7]  ( .D(n2403), .CLK(clk), .Q(\ram[209][7] ) );
  DFFNX1 \ram_reg[209][6]  ( .D(n2402), .CLK(clk), .Q(\ram[209][6] ) );
  DFFNX1 \ram_reg[209][5]  ( .D(n2401), .CLK(clk), .Q(\ram[209][5] ) );
  DFFNX1 \ram_reg[209][4]  ( .D(n2400), .CLK(clk), .Q(\ram[209][4] ) );
  DFFNX1 \ram_reg[209][3]  ( .D(n2399), .CLK(clk), .Q(\ram[209][3] ) );
  DFFNX1 \ram_reg[209][2]  ( .D(n2398), .CLK(clk), .Q(\ram[209][2] ) );
  DFFNX1 \ram_reg[209][1]  ( .D(n2397), .CLK(clk), .Q(\ram[209][1] ) );
  DFFNX1 \ram_reg[209][0]  ( .D(n2396), .CLK(clk), .Q(\ram[209][0] ) );
  DFFNX1 \ram_reg[210][7]  ( .D(n2395), .CLK(clk), .Q(\ram[210][7] ) );
  DFFNX1 \ram_reg[210][6]  ( .D(n2394), .CLK(clk), .Q(\ram[210][6] ) );
  DFFNX1 \ram_reg[210][5]  ( .D(n2393), .CLK(clk), .Q(\ram[210][5] ) );
  DFFNX1 \ram_reg[210][4]  ( .D(n2392), .CLK(clk), .Q(\ram[210][4] ) );
  DFFNX1 \ram_reg[210][3]  ( .D(n2391), .CLK(clk), .Q(\ram[210][3] ) );
  DFFNX1 \ram_reg[210][2]  ( .D(n2390), .CLK(clk), .Q(\ram[210][2] ) );
  DFFNX1 \ram_reg[210][1]  ( .D(n2389), .CLK(clk), .Q(\ram[210][1] ) );
  DFFNX1 \ram_reg[210][0]  ( .D(n2388), .CLK(clk), .Q(\ram[210][0] ) );
  DFFNX1 \ram_reg[211][7]  ( .D(n2387), .CLK(clk), .Q(\ram[211][7] ) );
  DFFNX1 \ram_reg[211][6]  ( .D(n2386), .CLK(clk), .Q(\ram[211][6] ) );
  DFFNX1 \ram_reg[211][5]  ( .D(n2385), .CLK(clk), .Q(\ram[211][5] ) );
  DFFNX1 \ram_reg[211][4]  ( .D(n2384), .CLK(clk), .Q(\ram[211][4] ) );
  DFFNX1 \ram_reg[211][3]  ( .D(n2383), .CLK(clk), .Q(\ram[211][3] ) );
  DFFNX1 \ram_reg[211][2]  ( .D(n2382), .CLK(clk), .Q(\ram[211][2] ) );
  DFFNX1 \ram_reg[211][1]  ( .D(n2381), .CLK(clk), .Q(\ram[211][1] ) );
  DFFNX1 \ram_reg[211][0]  ( .D(n2380), .CLK(clk), .Q(\ram[211][0] ) );
  DFFNX1 \ram_reg[212][7]  ( .D(n2379), .CLK(clk), .Q(\ram[212][7] ) );
  DFFNX1 \ram_reg[212][6]  ( .D(n2378), .CLK(clk), .Q(\ram[212][6] ) );
  DFFNX1 \ram_reg[212][5]  ( .D(n2377), .CLK(clk), .Q(\ram[212][5] ) );
  DFFNX1 \ram_reg[212][4]  ( .D(n2376), .CLK(clk), .Q(\ram[212][4] ) );
  DFFNX1 \ram_reg[212][3]  ( .D(n2375), .CLK(clk), .Q(\ram[212][3] ) );
  DFFNX1 \ram_reg[212][2]  ( .D(n2374), .CLK(clk), .Q(\ram[212][2] ) );
  DFFNX1 \ram_reg[212][1]  ( .D(n2373), .CLK(clk), .Q(\ram[212][1] ) );
  DFFNX1 \ram_reg[212][0]  ( .D(n2372), .CLK(clk), .Q(\ram[212][0] ) );
  DFFNX1 \ram_reg[213][7]  ( .D(n2371), .CLK(clk), .Q(\ram[213][7] ) );
  DFFNX1 \ram_reg[213][6]  ( .D(n2370), .CLK(clk), .Q(\ram[213][6] ) );
  DFFNX1 \ram_reg[213][5]  ( .D(n2369), .CLK(clk), .Q(\ram[213][5] ) );
  DFFNX1 \ram_reg[213][4]  ( .D(n2368), .CLK(clk), .Q(\ram[213][4] ) );
  DFFNX1 \ram_reg[213][3]  ( .D(n2367), .CLK(clk), .Q(\ram[213][3] ) );
  DFFNX1 \ram_reg[213][2]  ( .D(n2366), .CLK(clk), .Q(\ram[213][2] ) );
  DFFNX1 \ram_reg[213][1]  ( .D(n2365), .CLK(clk), .Q(\ram[213][1] ) );
  DFFNX1 \ram_reg[213][0]  ( .D(n2364), .CLK(clk), .Q(\ram[213][0] ) );
  DFFNX1 \ram_reg[214][7]  ( .D(n2363), .CLK(clk), .Q(\ram[214][7] ) );
  DFFNX1 \ram_reg[214][6]  ( .D(n2362), .CLK(clk), .Q(\ram[214][6] ) );
  DFFNX1 \ram_reg[214][5]  ( .D(n2361), .CLK(clk), .Q(\ram[214][5] ) );
  DFFNX1 \ram_reg[214][4]  ( .D(n2360), .CLK(clk), .Q(\ram[214][4] ) );
  DFFNX1 \ram_reg[214][3]  ( .D(n2359), .CLK(clk), .Q(\ram[214][3] ) );
  DFFNX1 \ram_reg[214][2]  ( .D(n2358), .CLK(clk), .Q(\ram[214][2] ) );
  DFFNX1 \ram_reg[214][1]  ( .D(n2357), .CLK(clk), .Q(\ram[214][1] ) );
  DFFNX1 \ram_reg[214][0]  ( .D(n2356), .CLK(clk), .Q(\ram[214][0] ) );
  DFFNX1 \ram_reg[215][7]  ( .D(n2355), .CLK(clk), .Q(\ram[215][7] ) );
  DFFNX1 \ram_reg[215][6]  ( .D(n2354), .CLK(clk), .Q(\ram[215][6] ) );
  DFFNX1 \ram_reg[215][5]  ( .D(n2353), .CLK(clk), .Q(\ram[215][5] ) );
  DFFNX1 \ram_reg[215][4]  ( .D(n2352), .CLK(clk), .Q(\ram[215][4] ) );
  DFFNX1 \ram_reg[215][3]  ( .D(n2351), .CLK(clk), .Q(\ram[215][3] ) );
  DFFNX1 \ram_reg[215][2]  ( .D(n2350), .CLK(clk), .Q(\ram[215][2] ) );
  DFFNX1 \ram_reg[215][1]  ( .D(n2349), .CLK(clk), .Q(\ram[215][1] ) );
  DFFNX1 \ram_reg[215][0]  ( .D(n2348), .CLK(clk), .Q(\ram[215][0] ) );
  DFFNX1 \ram_reg[216][7]  ( .D(n2347), .CLK(clk), .Q(\ram[216][7] ) );
  DFFNX1 \ram_reg[216][6]  ( .D(n2346), .CLK(clk), .Q(\ram[216][6] ) );
  DFFNX1 \ram_reg[216][5]  ( .D(n2345), .CLK(clk), .Q(\ram[216][5] ) );
  DFFNX1 \ram_reg[216][4]  ( .D(n2344), .CLK(clk), .Q(\ram[216][4] ) );
  DFFNX1 \ram_reg[216][3]  ( .D(n2343), .CLK(clk), .Q(\ram[216][3] ) );
  DFFNX1 \ram_reg[216][2]  ( .D(n2342), .CLK(clk), .Q(\ram[216][2] ) );
  DFFNX1 \ram_reg[216][1]  ( .D(n2341), .CLK(clk), .Q(\ram[216][1] ) );
  DFFNX1 \ram_reg[216][0]  ( .D(n2340), .CLK(clk), .Q(\ram[216][0] ) );
  DFFNX1 \ram_reg[217][7]  ( .D(n2339), .CLK(clk), .Q(\ram[217][7] ) );
  DFFNX1 \ram_reg[217][6]  ( .D(n2338), .CLK(clk), .Q(\ram[217][6] ) );
  DFFNX1 \ram_reg[217][5]  ( .D(n2337), .CLK(clk), .Q(\ram[217][5] ) );
  DFFNX1 \ram_reg[217][4]  ( .D(n2336), .CLK(clk), .Q(\ram[217][4] ) );
  DFFNX1 \ram_reg[217][3]  ( .D(n2335), .CLK(clk), .Q(\ram[217][3] ) );
  DFFNX1 \ram_reg[217][2]  ( .D(n2334), .CLK(clk), .Q(\ram[217][2] ) );
  DFFNX1 \ram_reg[217][1]  ( .D(n2333), .CLK(clk), .Q(\ram[217][1] ) );
  DFFNX1 \ram_reg[217][0]  ( .D(n2332), .CLK(clk), .Q(\ram[217][0] ) );
  DFFNX1 \ram_reg[218][7]  ( .D(n2331), .CLK(clk), .Q(\ram[218][7] ) );
  DFFNX1 \ram_reg[218][6]  ( .D(n2330), .CLK(clk), .Q(\ram[218][6] ) );
  DFFNX1 \ram_reg[218][5]  ( .D(n2329), .CLK(clk), .Q(\ram[218][5] ) );
  DFFNX1 \ram_reg[218][4]  ( .D(n2328), .CLK(clk), .Q(\ram[218][4] ) );
  DFFNX1 \ram_reg[218][3]  ( .D(n2327), .CLK(clk), .Q(\ram[218][3] ) );
  DFFNX1 \ram_reg[218][2]  ( .D(n2326), .CLK(clk), .Q(\ram[218][2] ) );
  DFFNX1 \ram_reg[218][1]  ( .D(n2325), .CLK(clk), .Q(\ram[218][1] ) );
  DFFNX1 \ram_reg[218][0]  ( .D(n2324), .CLK(clk), .Q(\ram[218][0] ) );
  DFFNX1 \ram_reg[219][7]  ( .D(n2323), .CLK(clk), .Q(\ram[219][7] ) );
  DFFNX1 \ram_reg[219][6]  ( .D(n2322), .CLK(clk), .Q(\ram[219][6] ) );
  DFFNX1 \ram_reg[219][5]  ( .D(n2321), .CLK(clk), .Q(\ram[219][5] ) );
  DFFNX1 \ram_reg[219][4]  ( .D(n2320), .CLK(clk), .Q(\ram[219][4] ) );
  DFFNX1 \ram_reg[219][3]  ( .D(n2319), .CLK(clk), .Q(\ram[219][3] ) );
  DFFNX1 \ram_reg[219][2]  ( .D(n2318), .CLK(clk), .Q(\ram[219][2] ) );
  DFFNX1 \ram_reg[219][1]  ( .D(n2317), .CLK(clk), .Q(\ram[219][1] ) );
  DFFNX1 \ram_reg[219][0]  ( .D(n2316), .CLK(clk), .Q(\ram[219][0] ) );
  DFFNX1 \ram_reg[220][7]  ( .D(n2315), .CLK(clk), .Q(\ram[220][7] ) );
  DFFNX1 \ram_reg[220][6]  ( .D(n2314), .CLK(clk), .Q(\ram[220][6] ) );
  DFFNX1 \ram_reg[220][5]  ( .D(n2313), .CLK(clk), .Q(\ram[220][5] ) );
  DFFNX1 \ram_reg[220][4]  ( .D(n2312), .CLK(clk), .Q(\ram[220][4] ) );
  DFFNX1 \ram_reg[220][3]  ( .D(n2311), .CLK(clk), .Q(\ram[220][3] ) );
  DFFNX1 \ram_reg[220][2]  ( .D(n2310), .CLK(clk), .Q(\ram[220][2] ) );
  DFFNX1 \ram_reg[220][1]  ( .D(n2309), .CLK(clk), .Q(\ram[220][1] ) );
  DFFNX1 \ram_reg[220][0]  ( .D(n2308), .CLK(clk), .Q(\ram[220][0] ) );
  DFFNX1 \ram_reg[221][7]  ( .D(n2307), .CLK(clk), .Q(\ram[221][7] ) );
  DFFNX1 \ram_reg[221][6]  ( .D(n2306), .CLK(clk), .Q(\ram[221][6] ) );
  DFFNX1 \ram_reg[221][5]  ( .D(n2305), .CLK(clk), .Q(\ram[221][5] ) );
  DFFNX1 \ram_reg[221][4]  ( .D(n2304), .CLK(clk), .Q(\ram[221][4] ) );
  DFFNX1 \ram_reg[221][3]  ( .D(n2303), .CLK(clk), .Q(\ram[221][3] ) );
  DFFNX1 \ram_reg[221][2]  ( .D(n2302), .CLK(clk), .Q(\ram[221][2] ) );
  DFFNX1 \ram_reg[221][1]  ( .D(n2301), .CLK(clk), .Q(\ram[221][1] ) );
  DFFNX1 \ram_reg[221][0]  ( .D(n2300), .CLK(clk), .Q(\ram[221][0] ) );
  DFFNX1 \ram_reg[222][7]  ( .D(n2299), .CLK(clk), .Q(\ram[222][7] ) );
  DFFNX1 \ram_reg[222][6]  ( .D(n2298), .CLK(clk), .Q(\ram[222][6] ) );
  DFFNX1 \ram_reg[222][5]  ( .D(n2297), .CLK(clk), .Q(\ram[222][5] ) );
  DFFNX1 \ram_reg[222][4]  ( .D(n2296), .CLK(clk), .Q(\ram[222][4] ) );
  DFFNX1 \ram_reg[222][3]  ( .D(n2295), .CLK(clk), .Q(\ram[222][3] ) );
  DFFNX1 \ram_reg[222][2]  ( .D(n2294), .CLK(clk), .Q(\ram[222][2] ) );
  DFFNX1 \ram_reg[222][1]  ( .D(n2293), .CLK(clk), .Q(\ram[222][1] ) );
  DFFNX1 \ram_reg[222][0]  ( .D(n2292), .CLK(clk), .Q(\ram[222][0] ) );
  DFFNX1 \ram_reg[223][7]  ( .D(n2291), .CLK(clk), .Q(\ram[223][7] ) );
  DFFNX1 \ram_reg[223][6]  ( .D(n2290), .CLK(clk), .Q(\ram[223][6] ) );
  DFFNX1 \ram_reg[223][5]  ( .D(n2289), .CLK(clk), .Q(\ram[223][5] ) );
  DFFNX1 \ram_reg[223][4]  ( .D(n2288), .CLK(clk), .Q(\ram[223][4] ) );
  DFFNX1 \ram_reg[223][3]  ( .D(n2287), .CLK(clk), .Q(\ram[223][3] ) );
  DFFNX1 \ram_reg[223][2]  ( .D(n2286), .CLK(clk), .Q(\ram[223][2] ) );
  DFFNX1 \ram_reg[223][1]  ( .D(n2285), .CLK(clk), .Q(\ram[223][1] ) );
  DFFNX1 \ram_reg[223][0]  ( .D(n2284), .CLK(clk), .Q(\ram[223][0] ) );
  DFFNX1 \ram_reg[224][7]  ( .D(n2283), .CLK(clk), .Q(\ram[224][7] ) );
  DFFNX1 \ram_reg[224][6]  ( .D(n2282), .CLK(clk), .Q(\ram[224][6] ) );
  DFFNX1 \ram_reg[224][5]  ( .D(n2281), .CLK(clk), .Q(\ram[224][5] ) );
  DFFNX1 \ram_reg[224][4]  ( .D(n2280), .CLK(clk), .Q(\ram[224][4] ) );
  DFFNX1 \ram_reg[224][3]  ( .D(n2279), .CLK(clk), .Q(\ram[224][3] ) );
  DFFNX1 \ram_reg[224][2]  ( .D(n2278), .CLK(clk), .Q(\ram[224][2] ) );
  DFFNX1 \ram_reg[224][1]  ( .D(n2277), .CLK(clk), .Q(\ram[224][1] ) );
  DFFNX1 \ram_reg[224][0]  ( .D(n2276), .CLK(clk), .Q(\ram[224][0] ) );
  DFFNX1 \ram_reg[225][7]  ( .D(n2275), .CLK(clk), .Q(\ram[225][7] ) );
  DFFNX1 \ram_reg[225][6]  ( .D(n2274), .CLK(clk), .Q(\ram[225][6] ) );
  DFFNX1 \ram_reg[225][5]  ( .D(n2273), .CLK(clk), .Q(\ram[225][5] ) );
  DFFNX1 \ram_reg[225][4]  ( .D(n2272), .CLK(clk), .Q(\ram[225][4] ) );
  DFFNX1 \ram_reg[225][3]  ( .D(n2271), .CLK(clk), .Q(\ram[225][3] ) );
  DFFNX1 \ram_reg[225][2]  ( .D(n2270), .CLK(clk), .Q(\ram[225][2] ) );
  DFFNX1 \ram_reg[225][1]  ( .D(n2269), .CLK(clk), .Q(\ram[225][1] ) );
  DFFNX1 \ram_reg[225][0]  ( .D(n2268), .CLK(clk), .Q(\ram[225][0] ) );
  DFFNX1 \ram_reg[226][7]  ( .D(n2267), .CLK(clk), .Q(\ram[226][7] ) );
  DFFNX1 \ram_reg[226][6]  ( .D(n2266), .CLK(clk), .Q(\ram[226][6] ) );
  DFFNX1 \ram_reg[226][5]  ( .D(n2265), .CLK(clk), .Q(\ram[226][5] ) );
  DFFNX1 \ram_reg[226][4]  ( .D(n2264), .CLK(clk), .Q(\ram[226][4] ) );
  DFFNX1 \ram_reg[226][3]  ( .D(n2263), .CLK(clk), .Q(\ram[226][3] ) );
  DFFNX1 \ram_reg[226][2]  ( .D(n2262), .CLK(clk), .Q(\ram[226][2] ) );
  DFFNX1 \ram_reg[226][1]  ( .D(n2261), .CLK(clk), .Q(\ram[226][1] ) );
  DFFNX1 \ram_reg[226][0]  ( .D(n2260), .CLK(clk), .Q(\ram[226][0] ) );
  DFFNX1 \ram_reg[227][7]  ( .D(n2259), .CLK(clk), .Q(\ram[227][7] ) );
  DFFNX1 \ram_reg[227][6]  ( .D(n2258), .CLK(clk), .Q(\ram[227][6] ) );
  DFFNX1 \ram_reg[227][5]  ( .D(n2257), .CLK(clk), .Q(\ram[227][5] ) );
  DFFNX1 \ram_reg[227][4]  ( .D(n2256), .CLK(clk), .Q(\ram[227][4] ) );
  DFFNX1 \ram_reg[227][3]  ( .D(n2255), .CLK(clk), .Q(\ram[227][3] ) );
  DFFNX1 \ram_reg[227][2]  ( .D(n2254), .CLK(clk), .Q(\ram[227][2] ) );
  DFFNX1 \ram_reg[227][1]  ( .D(n2253), .CLK(clk), .Q(\ram[227][1] ) );
  DFFNX1 \ram_reg[227][0]  ( .D(n2252), .CLK(clk), .Q(\ram[227][0] ) );
  DFFNX1 \ram_reg[228][7]  ( .D(n2251), .CLK(clk), .Q(\ram[228][7] ) );
  DFFNX1 \ram_reg[228][6]  ( .D(n2250), .CLK(clk), .Q(\ram[228][6] ) );
  DFFNX1 \ram_reg[228][5]  ( .D(n2249), .CLK(clk), .Q(\ram[228][5] ) );
  DFFNX1 \ram_reg[228][4]  ( .D(n2248), .CLK(clk), .Q(\ram[228][4] ) );
  DFFNX1 \ram_reg[228][3]  ( .D(n2247), .CLK(clk), .Q(\ram[228][3] ) );
  DFFNX1 \ram_reg[228][2]  ( .D(n2246), .CLK(clk), .Q(\ram[228][2] ) );
  DFFNX1 \ram_reg[228][1]  ( .D(n2245), .CLK(clk), .Q(\ram[228][1] ) );
  DFFNX1 \ram_reg[228][0]  ( .D(n2244), .CLK(clk), .Q(\ram[228][0] ) );
  DFFNX1 \ram_reg[229][7]  ( .D(n2243), .CLK(clk), .Q(\ram[229][7] ) );
  DFFNX1 \ram_reg[229][6]  ( .D(n2242), .CLK(clk), .Q(\ram[229][6] ) );
  DFFNX1 \ram_reg[229][5]  ( .D(n2241), .CLK(clk), .Q(\ram[229][5] ) );
  DFFNX1 \ram_reg[229][4]  ( .D(n2240), .CLK(clk), .Q(\ram[229][4] ) );
  DFFNX1 \ram_reg[229][3]  ( .D(n2239), .CLK(clk), .Q(\ram[229][3] ) );
  DFFNX1 \ram_reg[229][2]  ( .D(n2238), .CLK(clk), .Q(\ram[229][2] ) );
  DFFNX1 \ram_reg[229][1]  ( .D(n2237), .CLK(clk), .Q(\ram[229][1] ) );
  DFFNX1 \ram_reg[229][0]  ( .D(n2236), .CLK(clk), .Q(\ram[229][0] ) );
  DFFNX1 \ram_reg[230][7]  ( .D(n2235), .CLK(clk), .Q(\ram[230][7] ) );
  DFFNX1 \ram_reg[230][6]  ( .D(n2234), .CLK(clk), .Q(\ram[230][6] ) );
  DFFNX1 \ram_reg[230][5]  ( .D(n2233), .CLK(clk), .Q(\ram[230][5] ) );
  DFFNX1 \ram_reg[230][4]  ( .D(n2232), .CLK(clk), .Q(\ram[230][4] ) );
  DFFNX1 \ram_reg[230][3]  ( .D(n2231), .CLK(clk), .Q(\ram[230][3] ) );
  DFFNX1 \ram_reg[230][2]  ( .D(n2230), .CLK(clk), .Q(\ram[230][2] ) );
  DFFNX1 \ram_reg[230][1]  ( .D(n2229), .CLK(clk), .Q(\ram[230][1] ) );
  DFFNX1 \ram_reg[230][0]  ( .D(n2228), .CLK(clk), .Q(\ram[230][0] ) );
  DFFNX1 \ram_reg[231][7]  ( .D(n2227), .CLK(clk), .Q(\ram[231][7] ) );
  DFFNX1 \ram_reg[231][6]  ( .D(n2226), .CLK(clk), .Q(\ram[231][6] ) );
  DFFNX1 \ram_reg[231][5]  ( .D(n2225), .CLK(clk), .Q(\ram[231][5] ) );
  DFFNX1 \ram_reg[231][4]  ( .D(n2224), .CLK(clk), .Q(\ram[231][4] ) );
  DFFNX1 \ram_reg[231][3]  ( .D(n2223), .CLK(clk), .Q(\ram[231][3] ) );
  DFFNX1 \ram_reg[231][2]  ( .D(n2222), .CLK(clk), .Q(\ram[231][2] ) );
  DFFNX1 \ram_reg[231][1]  ( .D(n2221), .CLK(clk), .Q(\ram[231][1] ) );
  DFFNX1 \ram_reg[231][0]  ( .D(n2220), .CLK(clk), .Q(\ram[231][0] ) );
  DFFNX1 \ram_reg[232][7]  ( .D(n2219), .CLK(clk), .Q(\ram[232][7] ) );
  DFFNX1 \ram_reg[232][6]  ( .D(n2218), .CLK(clk), .Q(\ram[232][6] ) );
  DFFNX1 \ram_reg[232][5]  ( .D(n2217), .CLK(clk), .Q(\ram[232][5] ) );
  DFFNX1 \ram_reg[232][4]  ( .D(n2216), .CLK(clk), .Q(\ram[232][4] ) );
  DFFNX1 \ram_reg[232][3]  ( .D(n2215), .CLK(clk), .Q(\ram[232][3] ) );
  DFFNX1 \ram_reg[232][2]  ( .D(n2214), .CLK(clk), .Q(\ram[232][2] ) );
  DFFNX1 \ram_reg[232][1]  ( .D(n2213), .CLK(clk), .Q(\ram[232][1] ) );
  DFFNX1 \ram_reg[232][0]  ( .D(n2212), .CLK(clk), .Q(\ram[232][0] ) );
  DFFNX1 \ram_reg[233][7]  ( .D(n2211), .CLK(clk), .Q(\ram[233][7] ) );
  DFFNX1 \ram_reg[233][6]  ( .D(n2210), .CLK(clk), .Q(\ram[233][6] ) );
  DFFNX1 \ram_reg[233][5]  ( .D(n2209), .CLK(clk), .Q(\ram[233][5] ) );
  DFFNX1 \ram_reg[233][4]  ( .D(n2208), .CLK(clk), .Q(\ram[233][4] ) );
  DFFNX1 \ram_reg[233][3]  ( .D(n2207), .CLK(clk), .Q(\ram[233][3] ) );
  DFFNX1 \ram_reg[233][2]  ( .D(n2206), .CLK(clk), .Q(\ram[233][2] ) );
  DFFNX1 \ram_reg[233][1]  ( .D(n2205), .CLK(clk), .Q(\ram[233][1] ) );
  DFFNX1 \ram_reg[233][0]  ( .D(n2204), .CLK(clk), .Q(\ram[233][0] ) );
  DFFNX1 \ram_reg[234][7]  ( .D(n2203), .CLK(clk), .Q(\ram[234][7] ) );
  DFFNX1 \ram_reg[234][6]  ( .D(n2202), .CLK(clk), .Q(\ram[234][6] ) );
  DFFNX1 \ram_reg[234][5]  ( .D(n2201), .CLK(clk), .Q(\ram[234][5] ) );
  DFFNX1 \ram_reg[234][4]  ( .D(n2200), .CLK(clk), .Q(\ram[234][4] ) );
  DFFNX1 \ram_reg[234][3]  ( .D(n2199), .CLK(clk), .Q(\ram[234][3] ) );
  DFFNX1 \ram_reg[234][2]  ( .D(n2198), .CLK(clk), .Q(\ram[234][2] ) );
  DFFNX1 \ram_reg[234][1]  ( .D(n2197), .CLK(clk), .Q(\ram[234][1] ) );
  DFFNX1 \ram_reg[234][0]  ( .D(n2196), .CLK(clk), .Q(\ram[234][0] ) );
  DFFNX1 \ram_reg[235][7]  ( .D(n2195), .CLK(clk), .Q(\ram[235][7] ) );
  DFFNX1 \ram_reg[235][6]  ( .D(n2194), .CLK(clk), .Q(\ram[235][6] ) );
  DFFNX1 \ram_reg[235][5]  ( .D(n2193), .CLK(clk), .Q(\ram[235][5] ) );
  DFFNX1 \ram_reg[235][4]  ( .D(n2192), .CLK(clk), .Q(\ram[235][4] ) );
  DFFNX1 \ram_reg[235][3]  ( .D(n2191), .CLK(clk), .Q(\ram[235][3] ) );
  DFFNX1 \ram_reg[235][2]  ( .D(n2190), .CLK(clk), .Q(\ram[235][2] ) );
  DFFNX1 \ram_reg[235][1]  ( .D(n2189), .CLK(clk), .Q(\ram[235][1] ) );
  DFFNX1 \ram_reg[235][0]  ( .D(n2188), .CLK(clk), .Q(\ram[235][0] ) );
  DFFNX1 \ram_reg[236][7]  ( .D(n2187), .CLK(clk), .Q(\ram[236][7] ) );
  DFFNX1 \ram_reg[236][6]  ( .D(n2186), .CLK(clk), .Q(\ram[236][6] ) );
  DFFNX1 \ram_reg[236][5]  ( .D(n2185), .CLK(clk), .Q(\ram[236][5] ) );
  DFFNX1 \ram_reg[236][4]  ( .D(n2184), .CLK(clk), .Q(\ram[236][4] ) );
  DFFNX1 \ram_reg[236][3]  ( .D(n2183), .CLK(clk), .Q(\ram[236][3] ) );
  DFFNX1 \ram_reg[236][2]  ( .D(n2182), .CLK(clk), .Q(\ram[236][2] ) );
  DFFNX1 \ram_reg[236][1]  ( .D(n2181), .CLK(clk), .Q(\ram[236][1] ) );
  DFFNX1 \ram_reg[236][0]  ( .D(n2180), .CLK(clk), .Q(\ram[236][0] ) );
  DFFNX1 \ram_reg[237][7]  ( .D(n2179), .CLK(clk), .Q(\ram[237][7] ) );
  DFFNX1 \ram_reg[237][6]  ( .D(n2178), .CLK(clk), .Q(\ram[237][6] ) );
  DFFNX1 \ram_reg[237][5]  ( .D(n2177), .CLK(clk), .Q(\ram[237][5] ) );
  DFFNX1 \ram_reg[237][4]  ( .D(n2176), .CLK(clk), .Q(\ram[237][4] ) );
  DFFNX1 \ram_reg[237][3]  ( .D(n2175), .CLK(clk), .Q(\ram[237][3] ) );
  DFFNX1 \ram_reg[237][2]  ( .D(n2174), .CLK(clk), .Q(\ram[237][2] ) );
  DFFNX1 \ram_reg[237][1]  ( .D(n2173), .CLK(clk), .Q(\ram[237][1] ) );
  DFFNX1 \ram_reg[237][0]  ( .D(n2172), .CLK(clk), .Q(\ram[237][0] ) );
  DFFNX1 \ram_reg[238][7]  ( .D(n2171), .CLK(clk), .Q(\ram[238][7] ) );
  DFFNX1 \ram_reg[238][6]  ( .D(n2170), .CLK(clk), .Q(\ram[238][6] ) );
  DFFNX1 \ram_reg[238][5]  ( .D(n2169), .CLK(clk), .Q(\ram[238][5] ) );
  DFFNX1 \ram_reg[238][4]  ( .D(n2168), .CLK(clk), .Q(\ram[238][4] ) );
  DFFNX1 \ram_reg[238][3]  ( .D(n2167), .CLK(clk), .Q(\ram[238][3] ) );
  DFFNX1 \ram_reg[238][2]  ( .D(n2166), .CLK(clk), .Q(\ram[238][2] ) );
  DFFNX1 \ram_reg[238][1]  ( .D(n2165), .CLK(clk), .Q(\ram[238][1] ) );
  DFFNX1 \ram_reg[238][0]  ( .D(n2164), .CLK(clk), .Q(\ram[238][0] ) );
  DFFNX1 \ram_reg[239][7]  ( .D(n2163), .CLK(clk), .Q(\ram[239][7] ) );
  DFFNX1 \ram_reg[239][6]  ( .D(n2162), .CLK(clk), .Q(\ram[239][6] ) );
  DFFNX1 \ram_reg[239][5]  ( .D(n2161), .CLK(clk), .Q(\ram[239][5] ) );
  DFFNX1 \ram_reg[239][4]  ( .D(n2160), .CLK(clk), .Q(\ram[239][4] ) );
  DFFNX1 \ram_reg[239][3]  ( .D(n2159), .CLK(clk), .Q(\ram[239][3] ) );
  DFFNX1 \ram_reg[239][2]  ( .D(n2158), .CLK(clk), .Q(\ram[239][2] ) );
  DFFNX1 \ram_reg[239][1]  ( .D(n2157), .CLK(clk), .Q(\ram[239][1] ) );
  DFFNX1 \ram_reg[239][0]  ( .D(n2156), .CLK(clk), .Q(\ram[239][0] ) );
  DFFNX1 \ram_reg[240][7]  ( .D(n2155), .CLK(clk), .Q(\ram[240][7] ) );
  DFFNX1 \ram_reg[240][6]  ( .D(n2154), .CLK(clk), .Q(\ram[240][6] ) );
  DFFNX1 \ram_reg[240][5]  ( .D(n2153), .CLK(clk), .Q(\ram[240][5] ) );
  DFFNX1 \ram_reg[240][4]  ( .D(n2152), .CLK(clk), .Q(\ram[240][4] ) );
  DFFNX1 \ram_reg[240][3]  ( .D(n2151), .CLK(clk), .Q(\ram[240][3] ) );
  DFFNX1 \ram_reg[240][2]  ( .D(n2150), .CLK(clk), .Q(\ram[240][2] ) );
  DFFNX1 \ram_reg[240][1]  ( .D(n2149), .CLK(clk), .Q(\ram[240][1] ) );
  DFFNX1 \ram_reg[240][0]  ( .D(n2148), .CLK(clk), .Q(\ram[240][0] ) );
  DFFNX1 \ram_reg[241][7]  ( .D(n2147), .CLK(clk), .Q(\ram[241][7] ) );
  DFFNX1 \ram_reg[241][6]  ( .D(n2146), .CLK(clk), .Q(\ram[241][6] ) );
  DFFNX1 \ram_reg[241][5]  ( .D(n2145), .CLK(clk), .Q(\ram[241][5] ) );
  DFFNX1 \ram_reg[241][4]  ( .D(n2144), .CLK(clk), .Q(\ram[241][4] ) );
  DFFNX1 \ram_reg[241][3]  ( .D(n2143), .CLK(clk), .Q(\ram[241][3] ) );
  DFFNX1 \ram_reg[241][2]  ( .D(n2142), .CLK(clk), .Q(\ram[241][2] ) );
  DFFNX1 \ram_reg[241][1]  ( .D(n2141), .CLK(clk), .Q(\ram[241][1] ) );
  DFFNX1 \ram_reg[241][0]  ( .D(n2140), .CLK(clk), .Q(\ram[241][0] ) );
  DFFNX1 \ram_reg[242][7]  ( .D(n2139), .CLK(clk), .Q(\ram[242][7] ) );
  DFFNX1 \ram_reg[242][6]  ( .D(n2138), .CLK(clk), .Q(\ram[242][6] ) );
  DFFNX1 \ram_reg[242][5]  ( .D(n2137), .CLK(clk), .Q(\ram[242][5] ) );
  DFFNX1 \ram_reg[242][4]  ( .D(n2136), .CLK(clk), .Q(\ram[242][4] ) );
  DFFNX1 \ram_reg[242][3]  ( .D(n2135), .CLK(clk), .Q(\ram[242][3] ) );
  DFFNX1 \ram_reg[242][2]  ( .D(n2134), .CLK(clk), .Q(\ram[242][2] ) );
  DFFNX1 \ram_reg[242][1]  ( .D(n2133), .CLK(clk), .Q(\ram[242][1] ) );
  DFFNX1 \ram_reg[242][0]  ( .D(n2132), .CLK(clk), .Q(\ram[242][0] ) );
  DFFNX1 \ram_reg[243][7]  ( .D(n2131), .CLK(clk), .Q(\ram[243][7] ) );
  DFFNX1 \ram_reg[243][6]  ( .D(n2130), .CLK(clk), .Q(\ram[243][6] ) );
  DFFNX1 \ram_reg[243][5]  ( .D(n2129), .CLK(clk), .Q(\ram[243][5] ) );
  DFFNX1 \ram_reg[243][4]  ( .D(n2128), .CLK(clk), .Q(\ram[243][4] ) );
  DFFNX1 \ram_reg[243][3]  ( .D(n2127), .CLK(clk), .Q(\ram[243][3] ) );
  DFFNX1 \ram_reg[243][2]  ( .D(n2126), .CLK(clk), .Q(\ram[243][2] ) );
  DFFNX1 \ram_reg[243][1]  ( .D(n2125), .CLK(clk), .Q(\ram[243][1] ) );
  DFFNX1 \ram_reg[243][0]  ( .D(n2124), .CLK(clk), .Q(\ram[243][0] ) );
  DFFNX1 \ram_reg[244][7]  ( .D(n2123), .CLK(clk), .Q(\ram[244][7] ) );
  DFFNX1 \ram_reg[244][6]  ( .D(n2122), .CLK(clk), .Q(\ram[244][6] ) );
  DFFNX1 \ram_reg[244][5]  ( .D(n2121), .CLK(clk), .Q(\ram[244][5] ) );
  DFFNX1 \ram_reg[244][4]  ( .D(n2120), .CLK(clk), .Q(\ram[244][4] ) );
  DFFNX1 \ram_reg[244][3]  ( .D(n2119), .CLK(clk), .Q(\ram[244][3] ) );
  DFFNX1 \ram_reg[244][2]  ( .D(n2118), .CLK(clk), .Q(\ram[244][2] ) );
  DFFNX1 \ram_reg[244][1]  ( .D(n2117), .CLK(clk), .Q(\ram[244][1] ) );
  DFFNX1 \ram_reg[244][0]  ( .D(n2116), .CLK(clk), .Q(\ram[244][0] ) );
  DFFNX1 \ram_reg[245][7]  ( .D(n2115), .CLK(clk), .Q(\ram[245][7] ) );
  DFFNX1 \ram_reg[245][6]  ( .D(n2114), .CLK(clk), .Q(\ram[245][6] ) );
  DFFNX1 \ram_reg[245][5]  ( .D(n2113), .CLK(clk), .Q(\ram[245][5] ) );
  DFFNX1 \ram_reg[245][4]  ( .D(n2112), .CLK(clk), .Q(\ram[245][4] ) );
  DFFNX1 \ram_reg[245][3]  ( .D(n2111), .CLK(clk), .Q(\ram[245][3] ) );
  DFFNX1 \ram_reg[245][2]  ( .D(n2110), .CLK(clk), .Q(\ram[245][2] ) );
  DFFNX1 \ram_reg[245][1]  ( .D(n2109), .CLK(clk), .Q(\ram[245][1] ) );
  DFFNX1 \ram_reg[245][0]  ( .D(n2108), .CLK(clk), .Q(\ram[245][0] ) );
  DFFNX1 \ram_reg[246][7]  ( .D(n2107), .CLK(clk), .Q(\ram[246][7] ) );
  DFFNX1 \ram_reg[246][6]  ( .D(n2106), .CLK(clk), .Q(\ram[246][6] ) );
  DFFNX1 \ram_reg[246][5]  ( .D(n2105), .CLK(clk), .Q(\ram[246][5] ) );
  DFFNX1 \ram_reg[246][4]  ( .D(n2104), .CLK(clk), .Q(\ram[246][4] ) );
  DFFNX1 \ram_reg[246][3]  ( .D(n2103), .CLK(clk), .Q(\ram[246][3] ) );
  DFFNX1 \ram_reg[246][2]  ( .D(n2102), .CLK(clk), .Q(\ram[246][2] ) );
  DFFNX1 \ram_reg[246][1]  ( .D(n2101), .CLK(clk), .Q(\ram[246][1] ) );
  DFFNX1 \ram_reg[246][0]  ( .D(n2100), .CLK(clk), .Q(\ram[246][0] ) );
  DFFNX1 \ram_reg[247][7]  ( .D(n2099), .CLK(clk), .Q(\ram[247][7] ) );
  DFFNX1 \ram_reg[247][6]  ( .D(n2098), .CLK(clk), .Q(\ram[247][6] ) );
  DFFNX1 \ram_reg[247][5]  ( .D(n2097), .CLK(clk), .Q(\ram[247][5] ) );
  DFFNX1 \ram_reg[247][4]  ( .D(n2096), .CLK(clk), .Q(\ram[247][4] ) );
  DFFNX1 \ram_reg[247][3]  ( .D(n2095), .CLK(clk), .Q(\ram[247][3] ) );
  DFFNX1 \ram_reg[247][2]  ( .D(n2094), .CLK(clk), .Q(\ram[247][2] ) );
  DFFNX1 \ram_reg[247][1]  ( .D(n2093), .CLK(clk), .Q(\ram[247][1] ) );
  DFFNX1 \ram_reg[247][0]  ( .D(n2092), .CLK(clk), .Q(\ram[247][0] ) );
  DFFNX1 \ram_reg[248][7]  ( .D(n2091), .CLK(clk), .Q(\ram[248][7] ) );
  DFFNX1 \ram_reg[248][6]  ( .D(n2090), .CLK(clk), .Q(\ram[248][6] ) );
  DFFNX1 \ram_reg[248][5]  ( .D(n2089), .CLK(clk), .Q(\ram[248][5] ) );
  DFFNX1 \ram_reg[248][4]  ( .D(n2088), .CLK(clk), .Q(\ram[248][4] ) );
  DFFNX1 \ram_reg[248][3]  ( .D(n2087), .CLK(clk), .Q(\ram[248][3] ) );
  DFFNX1 \ram_reg[248][2]  ( .D(n2086), .CLK(clk), .Q(\ram[248][2] ) );
  DFFNX1 \ram_reg[248][1]  ( .D(n2085), .CLK(clk), .Q(\ram[248][1] ) );
  DFFNX1 \ram_reg[248][0]  ( .D(n2084), .CLK(clk), .Q(\ram[248][0] ) );
  DFFNX1 \ram_reg[249][7]  ( .D(n2083), .CLK(clk), .Q(\ram[249][7] ) );
  DFFNX1 \ram_reg[249][6]  ( .D(n2082), .CLK(clk), .Q(\ram[249][6] ) );
  DFFNX1 \ram_reg[249][5]  ( .D(n2081), .CLK(clk), .Q(\ram[249][5] ) );
  DFFNX1 \ram_reg[249][4]  ( .D(n2080), .CLK(clk), .Q(\ram[249][4] ) );
  DFFNX1 \ram_reg[249][3]  ( .D(n2079), .CLK(clk), .Q(\ram[249][3] ) );
  DFFNX1 \ram_reg[249][2]  ( .D(n2078), .CLK(clk), .Q(\ram[249][2] ) );
  DFFNX1 \ram_reg[249][1]  ( .D(n2077), .CLK(clk), .Q(\ram[249][1] ) );
  DFFNX1 \ram_reg[249][0]  ( .D(n2076), .CLK(clk), .Q(\ram[249][0] ) );
  DFFNX1 \ram_reg[250][7]  ( .D(n2075), .CLK(clk), .Q(\ram[250][7] ) );
  DFFNX1 \ram_reg[250][6]  ( .D(n2074), .CLK(clk), .Q(\ram[250][6] ) );
  DFFNX1 \ram_reg[250][5]  ( .D(n2073), .CLK(clk), .Q(\ram[250][5] ) );
  DFFNX1 \ram_reg[250][4]  ( .D(n2072), .CLK(clk), .Q(\ram[250][4] ) );
  DFFNX1 \ram_reg[250][3]  ( .D(n2071), .CLK(clk), .Q(\ram[250][3] ) );
  DFFNX1 \ram_reg[250][2]  ( .D(n2070), .CLK(clk), .Q(\ram[250][2] ) );
  DFFNX1 \ram_reg[250][1]  ( .D(n2069), .CLK(clk), .Q(\ram[250][1] ) );
  DFFNX1 \ram_reg[250][0]  ( .D(n2068), .CLK(clk), .Q(\ram[250][0] ) );
  DFFNX1 \ram_reg[251][7]  ( .D(n2067), .CLK(clk), .Q(\ram[251][7] ) );
  DFFNX1 \ram_reg[251][6]  ( .D(n2066), .CLK(clk), .Q(\ram[251][6] ) );
  DFFNX1 \ram_reg[251][5]  ( .D(n2065), .CLK(clk), .Q(\ram[251][5] ) );
  DFFNX1 \ram_reg[251][4]  ( .D(n2064), .CLK(clk), .Q(\ram[251][4] ) );
  DFFNX1 \ram_reg[251][3]  ( .D(n2063), .CLK(clk), .Q(\ram[251][3] ) );
  DFFNX1 \ram_reg[251][2]  ( .D(n2062), .CLK(clk), .Q(\ram[251][2] ) );
  DFFNX1 \ram_reg[251][1]  ( .D(n2061), .CLK(clk), .Q(\ram[251][1] ) );
  DFFNX1 \ram_reg[251][0]  ( .D(n2060), .CLK(clk), .Q(\ram[251][0] ) );
  DFFNX1 \ram_reg[252][7]  ( .D(n2059), .CLK(clk), .Q(\ram[252][7] ) );
  DFFNX1 \ram_reg[252][6]  ( .D(n2058), .CLK(clk), .Q(\ram[252][6] ) );
  DFFNX1 \ram_reg[252][5]  ( .D(n2057), .CLK(clk), .Q(\ram[252][5] ) );
  DFFNX1 \ram_reg[252][4]  ( .D(n2056), .CLK(clk), .Q(\ram[252][4] ) );
  DFFNX1 \ram_reg[252][3]  ( .D(n2055), .CLK(clk), .Q(\ram[252][3] ) );
  DFFNX1 \ram_reg[252][2]  ( .D(n2054), .CLK(clk), .Q(\ram[252][2] ) );
  DFFNX1 \ram_reg[252][1]  ( .D(n2053), .CLK(clk), .Q(\ram[252][1] ) );
  DFFNX1 \ram_reg[252][0]  ( .D(n2052), .CLK(clk), .Q(\ram[252][0] ) );
  DFFNX1 \ram_reg[253][7]  ( .D(n2051), .CLK(clk), .Q(\ram[253][7] ) );
  DFFNX1 \ram_reg[253][6]  ( .D(n2050), .CLK(clk), .Q(\ram[253][6] ) );
  DFFNX1 \ram_reg[253][5]  ( .D(n2049), .CLK(clk), .Q(\ram[253][5] ) );
  DFFNX1 \ram_reg[253][4]  ( .D(n2048), .CLK(clk), .Q(\ram[253][4] ) );
  DFFNX1 \ram_reg[253][3]  ( .D(n2047), .CLK(clk), .Q(\ram[253][3] ) );
  DFFNX1 \ram_reg[253][2]  ( .D(n2046), .CLK(clk), .Q(\ram[253][2] ) );
  DFFNX1 \ram_reg[253][1]  ( .D(n2045), .CLK(clk), .Q(\ram[253][1] ) );
  DFFNX1 \ram_reg[253][0]  ( .D(n2044), .CLK(clk), .Q(\ram[253][0] ) );
  DFFNX1 \ram_reg[254][7]  ( .D(n2043), .CLK(clk), .Q(\ram[254][7] ) );
  DFFNX1 \ram_reg[254][6]  ( .D(n2042), .CLK(clk), .Q(\ram[254][6] ) );
  DFFNX1 \ram_reg[254][5]  ( .D(n2041), .CLK(clk), .Q(\ram[254][5] ) );
  DFFNX1 \ram_reg[254][4]  ( .D(n2040), .CLK(clk), .Q(\ram[254][4] ) );
  DFFNX1 \ram_reg[254][3]  ( .D(n2039), .CLK(clk), .Q(\ram[254][3] ) );
  DFFNX1 \ram_reg[254][2]  ( .D(n2038), .CLK(clk), .Q(\ram[254][2] ) );
  DFFNX1 \ram_reg[254][1]  ( .D(n2037), .CLK(clk), .Q(\ram[254][1] ) );
  DFFNX1 \ram_reg[254][0]  ( .D(n2036), .CLK(clk), .Q(\ram[254][0] ) );
  DFFNX1 \ram_reg[255][7]  ( .D(n2035), .CLK(clk), .Q(\ram[255][7] ) );
  DFFNX1 \ram_reg[255][6]  ( .D(n2034), .CLK(clk), .Q(\ram[255][6] ) );
  DFFNX1 \ram_reg[255][5]  ( .D(n2033), .CLK(clk), .Q(\ram[255][5] ) );
  DFFNX1 \ram_reg[255][4]  ( .D(n2032), .CLK(clk), .Q(\ram[255][4] ) );
  DFFNX1 \ram_reg[255][3]  ( .D(n2031), .CLK(clk), .Q(\ram[255][3] ) );
  DFFNX1 \ram_reg[255][2]  ( .D(n2030), .CLK(clk), .Q(\ram[255][2] ) );
  DFFNX1 \ram_reg[255][1]  ( .D(n2029), .CLK(clk), .Q(\ram[255][1] ) );
  DFFNX1 \ram_reg[255][0]  ( .D(n2028), .CLK(clk), .Q(\ram[255][0] ) );
  DFFNX1 \dataout_reg[7]  ( .D(n2027), .CLK(clk), .Q(dataout[7]) );
  DFFNX1 \dataout_reg[6]  ( .D(n2026), .CLK(clk), .Q(dataout[6]) );
  DFFNX1 \dataout_reg[5]  ( .D(n2025), .CLK(clk), .Q(dataout[5]) );
  DFFNX1 \dataout_reg[4]  ( .D(n2024), .CLK(clk), .Q(dataout[4]) );
  DFFNX1 \dataout_reg[3]  ( .D(n2023), .CLK(clk), .Q(dataout[3]) );
  DFFNX1 \dataout_reg[2]  ( .D(n2022), .CLK(clk), .Q(dataout[2]) );
  DFFNX1 \dataout_reg[1]  ( .D(n2021), .CLK(clk), .Q(dataout[1]) );
  DFFNX1 \dataout_reg[0]  ( .D(n2020), .CLK(clk), .Q(dataout[0]) );
  DFFNX1 MFC_reg ( .D(n4174), .CLK(clk), .Q(MFC) );
  AO22X1 U3 ( .IN1(\ram[255][0] ), .IN2(n1), .IN3(datain[0]), .IN4(n387), .Q(
        n2028) );
  AO22X1 U4 ( .IN1(\ram[255][1] ), .IN2(n1), .IN3(datain[1]), .IN4(n387), .Q(
        n2029) );
  AO22X1 U5 ( .IN1(\ram[255][2] ), .IN2(n1), .IN3(datain[2]), .IN4(n387), .Q(
        n2030) );
  AO22X1 U6 ( .IN1(\ram[255][3] ), .IN2(n1), .IN3(datain[3]), .IN4(n387), .Q(
        n2031) );
  AO22X1 U7 ( .IN1(\ram[255][4] ), .IN2(n1), .IN3(datain[4]), .IN4(n387), .Q(
        n2032) );
  AO22X1 U8 ( .IN1(\ram[255][5] ), .IN2(n1), .IN3(datain[5]), .IN4(n387), .Q(
        n2033) );
  AO22X1 U9 ( .IN1(\ram[255][6] ), .IN2(n1), .IN3(datain[6]), .IN4(n387), .Q(
        n2034) );
  AO22X1 U10 ( .IN1(\ram[255][7] ), .IN2(n1), .IN3(datain[7]), .IN4(n387), .Q(
        n2035) );
  AO22X1 U13 ( .IN1(\ram[254][0] ), .IN2(n5), .IN3(n4087), .IN4(n57), .Q(n2036) );
  AO22X1 U14 ( .IN1(\ram[254][1] ), .IN2(n5), .IN3(n4087), .IN4(n90), .Q(n2037) );
  AO22X1 U15 ( .IN1(\ram[254][2] ), .IN2(n5), .IN3(n4087), .IN4(n123), .Q(
        n2038) );
  AO22X1 U16 ( .IN1(\ram[254][3] ), .IN2(n5), .IN3(n4087), .IN4(n156), .Q(
        n2039) );
  AO22X1 U17 ( .IN1(\ram[254][4] ), .IN2(n5), .IN3(n4087), .IN4(n189), .Q(
        n2040) );
  AO22X1 U18 ( .IN1(\ram[254][5] ), .IN2(n5), .IN3(n4087), .IN4(n222), .Q(
        n2041) );
  AO22X1 U19 ( .IN1(\ram[254][6] ), .IN2(n5), .IN3(n4087), .IN4(n255), .Q(
        n2042) );
  AO22X1 U20 ( .IN1(\ram[254][7] ), .IN2(n5), .IN3(n4087), .IN4(n288), .Q(
        n2043) );
  AO22X1 U23 ( .IN1(\ram[253][0] ), .IN2(n8), .IN3(n444), .IN4(n54), .Q(n2044)
         );
  AO22X1 U24 ( .IN1(\ram[253][1] ), .IN2(n8), .IN3(n444), .IN4(n87), .Q(n2045)
         );
  AO22X1 U25 ( .IN1(\ram[253][2] ), .IN2(n8), .IN3(n444), .IN4(n120), .Q(n2046) );
  AO22X1 U26 ( .IN1(\ram[253][3] ), .IN2(n8), .IN3(n444), .IN4(n153), .Q(n2047) );
  AO22X1 U27 ( .IN1(\ram[253][4] ), .IN2(n8), .IN3(n444), .IN4(n186), .Q(n2048) );
  AO22X1 U28 ( .IN1(\ram[253][5] ), .IN2(n8), .IN3(n444), .IN4(n219), .Q(n2049) );
  AO22X1 U29 ( .IN1(\ram[253][6] ), .IN2(n8), .IN3(n444), .IN4(n252), .Q(n2050) );
  AO22X1 U30 ( .IN1(\ram[253][7] ), .IN2(n8), .IN3(n444), .IN4(n285), .Q(n2051) );
  AO22X1 U33 ( .IN1(\ram[252][0] ), .IN2(n11), .IN3(n2006), .IN4(n60), .Q(
        n2052) );
  AO22X1 U34 ( .IN1(\ram[252][1] ), .IN2(n11), .IN3(n2006), .IN4(n93), .Q(
        n2053) );
  AO22X1 U35 ( .IN1(\ram[252][2] ), .IN2(n11), .IN3(n2006), .IN4(n126), .Q(
        n2054) );
  AO22X1 U36 ( .IN1(\ram[252][3] ), .IN2(n11), .IN3(n2006), .IN4(n159), .Q(
        n2055) );
  AO22X1 U37 ( .IN1(\ram[252][4] ), .IN2(n11), .IN3(n2006), .IN4(n192), .Q(
        n2056) );
  AO22X1 U38 ( .IN1(\ram[252][5] ), .IN2(n11), .IN3(n2006), .IN4(n225), .Q(
        n2057) );
  AO22X1 U39 ( .IN1(\ram[252][6] ), .IN2(n11), .IN3(n2006), .IN4(n258), .Q(
        n2058) );
  AO22X1 U40 ( .IN1(\ram[252][7] ), .IN2(n11), .IN3(n2006), .IN4(n291), .Q(
        n2059) );
  AO22X1 U43 ( .IN1(\ram[251][0] ), .IN2(n14), .IN3(n345), .IN4(n51), .Q(n2060) );
  AO22X1 U44 ( .IN1(\ram[251][1] ), .IN2(n14), .IN3(n345), .IN4(n84), .Q(n2061) );
  AO22X1 U45 ( .IN1(\ram[251][2] ), .IN2(n14), .IN3(n345), .IN4(n117), .Q(
        n2062) );
  AO22X1 U46 ( .IN1(\ram[251][3] ), .IN2(n14), .IN3(n345), .IN4(n150), .Q(
        n2063) );
  AO22X1 U47 ( .IN1(\ram[251][4] ), .IN2(n14), .IN3(n345), .IN4(n183), .Q(
        n2064) );
  AO22X1 U48 ( .IN1(\ram[251][5] ), .IN2(n14), .IN3(n345), .IN4(n216), .Q(
        n2065) );
  AO22X1 U49 ( .IN1(\ram[251][6] ), .IN2(n14), .IN3(n345), .IN4(n249), .Q(
        n2066) );
  AO22X1 U50 ( .IN1(\ram[251][7] ), .IN2(n14), .IN3(n345), .IN4(n282), .Q(
        n2067) );
  AO22X1 U53 ( .IN1(\ram[250][0] ), .IN2(n17), .IN3(n2007), .IN4(n48), .Q(
        n2068) );
  AO22X1 U54 ( .IN1(\ram[250][1] ), .IN2(n17), .IN3(n2007), .IN4(n81), .Q(
        n2069) );
  AO22X1 U55 ( .IN1(\ram[250][2] ), .IN2(n17), .IN3(n2007), .IN4(n114), .Q(
        n2070) );
  AO22X1 U56 ( .IN1(\ram[250][3] ), .IN2(n17), .IN3(n2007), .IN4(n147), .Q(
        n2071) );
  AO22X1 U57 ( .IN1(\ram[250][4] ), .IN2(n17), .IN3(n2007), .IN4(n180), .Q(
        n2072) );
  AO22X1 U58 ( .IN1(\ram[250][5] ), .IN2(n17), .IN3(n2007), .IN4(n213), .Q(
        n2073) );
  AO22X1 U59 ( .IN1(\ram[250][6] ), .IN2(n17), .IN3(n2007), .IN4(n246), .Q(
        n2074) );
  AO22X1 U60 ( .IN1(\ram[250][7] ), .IN2(n17), .IN3(n2007), .IN4(n279), .Q(
        n2075) );
  AO22X1 U63 ( .IN1(\ram[249][0] ), .IN2(n20), .IN3(n396), .IN4(n45), .Q(n2076) );
  AO22X1 U64 ( .IN1(\ram[249][1] ), .IN2(n20), .IN3(n396), .IN4(n78), .Q(n2077) );
  AO22X1 U65 ( .IN1(\ram[249][2] ), .IN2(n20), .IN3(n396), .IN4(n111), .Q(
        n2078) );
  AO22X1 U66 ( .IN1(\ram[249][3] ), .IN2(n20), .IN3(n396), .IN4(n144), .Q(
        n2079) );
  AO22X1 U67 ( .IN1(\ram[249][4] ), .IN2(n20), .IN3(n396), .IN4(n177), .Q(
        n2080) );
  AO22X1 U68 ( .IN1(\ram[249][5] ), .IN2(n20), .IN3(n396), .IN4(n210), .Q(
        n2081) );
  AO22X1 U69 ( .IN1(\ram[249][6] ), .IN2(n20), .IN3(n396), .IN4(n243), .Q(
        n2082) );
  AO22X1 U70 ( .IN1(\ram[249][7] ), .IN2(n20), .IN3(n396), .IN4(n276), .Q(
        n2083) );
  AO22X1 U73 ( .IN1(\ram[248][0] ), .IN2(n23), .IN3(n717), .IN4(n42), .Q(n2084) );
  AO22X1 U74 ( .IN1(\ram[248][1] ), .IN2(n23), .IN3(n717), .IN4(n75), .Q(n2085) );
  AO22X1 U75 ( .IN1(\ram[248][2] ), .IN2(n23), .IN3(n717), .IN4(n108), .Q(
        n2086) );
  AO22X1 U76 ( .IN1(\ram[248][3] ), .IN2(n23), .IN3(n717), .IN4(n141), .Q(
        n2087) );
  AO22X1 U77 ( .IN1(\ram[248][4] ), .IN2(n23), .IN3(n717), .IN4(n174), .Q(
        n2088) );
  AO22X1 U78 ( .IN1(\ram[248][5] ), .IN2(n23), .IN3(n717), .IN4(n207), .Q(
        n2089) );
  AO22X1 U79 ( .IN1(\ram[248][6] ), .IN2(n23), .IN3(n717), .IN4(n240), .Q(
        n2090) );
  AO22X1 U80 ( .IN1(\ram[248][7] ), .IN2(n23), .IN3(n717), .IN4(n273), .Q(
        n2091) );
  AO22X1 U83 ( .IN1(\ram[247][0] ), .IN2(n26), .IN3(n570), .IN4(n39), .Q(n2092) );
  AO22X1 U84 ( .IN1(\ram[247][1] ), .IN2(n26), .IN3(n570), .IN4(n72), .Q(n2093) );
  AO22X1 U85 ( .IN1(\ram[247][2] ), .IN2(n26), .IN3(n570), .IN4(n105), .Q(
        n2094) );
  AO22X1 U86 ( .IN1(\ram[247][3] ), .IN2(n26), .IN3(n570), .IN4(n138), .Q(
        n2095) );
  AO22X1 U87 ( .IN1(\ram[247][4] ), .IN2(n26), .IN3(n570), .IN4(n171), .Q(
        n2096) );
  AO22X1 U88 ( .IN1(\ram[247][5] ), .IN2(n26), .IN3(n570), .IN4(n204), .Q(
        n2097) );
  AO22X1 U89 ( .IN1(\ram[247][6] ), .IN2(n26), .IN3(n570), .IN4(n237), .Q(
        n2098) );
  AO22X1 U90 ( .IN1(\ram[247][7] ), .IN2(n26), .IN3(n570), .IN4(n270), .Q(
        n2099) );
  AO22X1 U93 ( .IN1(\ram[246][0] ), .IN2(n29), .IN3(n4161), .IN4(n36), .Q(
        n2100) );
  AO22X1 U94 ( .IN1(\ram[246][1] ), .IN2(n29), .IN3(n4161), .IN4(n69), .Q(
        n2101) );
  AO22X1 U95 ( .IN1(\ram[246][2] ), .IN2(n29), .IN3(n4161), .IN4(n102), .Q(
        n2102) );
  AO22X1 U96 ( .IN1(\ram[246][3] ), .IN2(n29), .IN3(n4161), .IN4(n135), .Q(
        n2103) );
  AO22X1 U97 ( .IN1(\ram[246][4] ), .IN2(n29), .IN3(n4161), .IN4(n168), .Q(
        n2104) );
  AO22X1 U98 ( .IN1(\ram[246][5] ), .IN2(n29), .IN3(n4161), .IN4(n201), .Q(
        n2105) );
  AO22X1 U99 ( .IN1(\ram[246][6] ), .IN2(n29), .IN3(n4161), .IN4(n234), .Q(
        n2106) );
  AO22X1 U100 ( .IN1(\ram[246][7] ), .IN2(n29), .IN3(n4161), .IN4(n267), .Q(
        n2107) );
  AO22X1 U103 ( .IN1(\ram[245][0] ), .IN2(n32), .IN3(n666), .IN4(datain[0]), 
        .Q(n2108) );
  AO22X1 U104 ( .IN1(\ram[245][1] ), .IN2(n32), .IN3(n666), .IN4(datain[1]), 
        .Q(n2109) );
  AO22X1 U105 ( .IN1(\ram[245][2] ), .IN2(n32), .IN3(n666), .IN4(datain[2]), 
        .Q(n2110) );
  AO22X1 U106 ( .IN1(\ram[245][3] ), .IN2(n32), .IN3(n666), .IN4(datain[3]), 
        .Q(n2111) );
  AO22X1 U107 ( .IN1(\ram[245][4] ), .IN2(n32), .IN3(n666), .IN4(datain[4]), 
        .Q(n2112) );
  AO22X1 U108 ( .IN1(\ram[245][5] ), .IN2(n32), .IN3(n666), .IN4(datain[5]), 
        .Q(n2113) );
  AO22X1 U109 ( .IN1(\ram[245][6] ), .IN2(n32), .IN3(n666), .IN4(datain[6]), 
        .Q(n2114) );
  AO22X1 U110 ( .IN1(\ram[245][7] ), .IN2(n32), .IN3(n666), .IN4(datain[7]), 
        .Q(n2115) );
  AO22X1 U113 ( .IN1(\ram[244][0] ), .IN2(n35), .IN3(n4113), .IN4(datain[0]), 
        .Q(n2116) );
  AO22X1 U114 ( .IN1(\ram[244][1] ), .IN2(n35), .IN3(n4113), .IN4(datain[1]), 
        .Q(n2117) );
  AO22X1 U115 ( .IN1(\ram[244][2] ), .IN2(n35), .IN3(n4113), .IN4(datain[2]), 
        .Q(n2118) );
  AO22X1 U116 ( .IN1(\ram[244][3] ), .IN2(n35), .IN3(n4113), .IN4(datain[3]), 
        .Q(n2119) );
  AO22X1 U117 ( .IN1(\ram[244][4] ), .IN2(n35), .IN3(n4113), .IN4(datain[4]), 
        .Q(n2120) );
  AO22X1 U118 ( .IN1(\ram[244][5] ), .IN2(n35), .IN3(n4113), .IN4(datain[5]), 
        .Q(n2121) );
  AO22X1 U119 ( .IN1(\ram[244][6] ), .IN2(n35), .IN3(n4113), .IN4(datain[6]), 
        .Q(n2122) );
  AO22X1 U120 ( .IN1(\ram[244][7] ), .IN2(n35), .IN3(n4113), .IN4(datain[7]), 
        .Q(n2123) );
  AO22X1 U123 ( .IN1(\ram[243][0] ), .IN2(n38), .IN3(n522), .IN4(datain[0]), 
        .Q(n2124) );
  AO22X1 U124 ( .IN1(\ram[243][1] ), .IN2(n38), .IN3(n522), .IN4(datain[1]), 
        .Q(n2125) );
  AO22X1 U125 ( .IN1(\ram[243][2] ), .IN2(n38), .IN3(n522), .IN4(datain[2]), 
        .Q(n2126) );
  AO22X1 U126 ( .IN1(\ram[243][3] ), .IN2(n38), .IN3(n522), .IN4(datain[3]), 
        .Q(n2127) );
  AO22X1 U127 ( .IN1(\ram[243][4] ), .IN2(n38), .IN3(n522), .IN4(datain[4]), 
        .Q(n2128) );
  AO22X1 U128 ( .IN1(\ram[243][5] ), .IN2(n38), .IN3(n522), .IN4(datain[5]), 
        .Q(n2129) );
  AO22X1 U129 ( .IN1(\ram[243][6] ), .IN2(n38), .IN3(n522), .IN4(datain[6]), 
        .Q(n2130) );
  AO22X1 U130 ( .IN1(\ram[243][7] ), .IN2(n38), .IN3(n522), .IN4(datain[7]), 
        .Q(n2131) );
  AO22X1 U133 ( .IN1(\ram[242][0] ), .IN2(n41), .IN3(n4144), .IN4(datain[0]), 
        .Q(n2132) );
  AO22X1 U134 ( .IN1(\ram[242][1] ), .IN2(n41), .IN3(n4144), .IN4(datain[1]), 
        .Q(n2133) );
  AO22X1 U135 ( .IN1(\ram[242][2] ), .IN2(n41), .IN3(n4144), .IN4(datain[2]), 
        .Q(n2134) );
  AO22X1 U136 ( .IN1(\ram[242][3] ), .IN2(n41), .IN3(n4144), .IN4(datain[3]), 
        .Q(n2135) );
  AO22X1 U137 ( .IN1(\ram[242][4] ), .IN2(n41), .IN3(n4144), .IN4(datain[4]), 
        .Q(n2136) );
  AO22X1 U138 ( .IN1(\ram[242][5] ), .IN2(n41), .IN3(n4144), .IN4(datain[5]), 
        .Q(n2137) );
  AO22X1 U139 ( .IN1(\ram[242][6] ), .IN2(n41), .IN3(n4144), .IN4(datain[6]), 
        .Q(n2138) );
  AO22X1 U140 ( .IN1(\ram[242][7] ), .IN2(n41), .IN3(n4144), .IN4(datain[7]), 
        .Q(n2139) );
  AO22X1 U143 ( .IN1(\ram[241][0] ), .IN2(n44), .IN3(n618), .IN4(datain[0]), 
        .Q(n2140) );
  AO22X1 U144 ( .IN1(\ram[241][1] ), .IN2(n44), .IN3(n618), .IN4(datain[1]), 
        .Q(n2141) );
  AO22X1 U145 ( .IN1(\ram[241][2] ), .IN2(n44), .IN3(n618), .IN4(datain[2]), 
        .Q(n2142) );
  AO22X1 U146 ( .IN1(\ram[241][3] ), .IN2(n44), .IN3(n618), .IN4(datain[3]), 
        .Q(n2143) );
  AO22X1 U147 ( .IN1(\ram[241][4] ), .IN2(n44), .IN3(n618), .IN4(datain[4]), 
        .Q(n2144) );
  AO22X1 U148 ( .IN1(\ram[241][5] ), .IN2(n44), .IN3(n618), .IN4(datain[5]), 
        .Q(n2145) );
  AO22X1 U149 ( .IN1(\ram[241][6] ), .IN2(n44), .IN3(n618), .IN4(datain[6]), 
        .Q(n2146) );
  AO22X1 U150 ( .IN1(\ram[241][7] ), .IN2(n44), .IN3(n618), .IN4(datain[7]), 
        .Q(n2147) );
  AO22X1 U153 ( .IN1(\ram[240][0] ), .IN2(n47), .IN3(n4133), .IN4(datain[0]), 
        .Q(n2148) );
  AO22X1 U154 ( .IN1(\ram[240][1] ), .IN2(n47), .IN3(n4133), .IN4(datain[1]), 
        .Q(n2149) );
  AO22X1 U155 ( .IN1(\ram[240][2] ), .IN2(n47), .IN3(n4133), .IN4(datain[2]), 
        .Q(n2150) );
  AO22X1 U156 ( .IN1(\ram[240][3] ), .IN2(n47), .IN3(n4133), .IN4(datain[3]), 
        .Q(n2151) );
  AO22X1 U157 ( .IN1(\ram[240][4] ), .IN2(n47), .IN3(n4133), .IN4(datain[4]), 
        .Q(n2152) );
  AO22X1 U158 ( .IN1(\ram[240][5] ), .IN2(n47), .IN3(n4133), .IN4(datain[5]), 
        .Q(n2153) );
  AO22X1 U159 ( .IN1(\ram[240][6] ), .IN2(n47), .IN3(n4133), .IN4(datain[6]), 
        .Q(n2154) );
  AO22X1 U160 ( .IN1(\ram[240][7] ), .IN2(n47), .IN3(n4133), .IN4(datain[7]), 
        .Q(n2155) );
  AO22X1 U163 ( .IN1(\ram[239][0] ), .IN2(n50), .IN3(n390), .IN4(datain[0]), 
        .Q(n2156) );
  AO22X1 U164 ( .IN1(\ram[239][1] ), .IN2(n50), .IN3(n390), .IN4(datain[1]), 
        .Q(n2157) );
  AO22X1 U165 ( .IN1(\ram[239][2] ), .IN2(n50), .IN3(n390), .IN4(datain[2]), 
        .Q(n2158) );
  AO22X1 U166 ( .IN1(\ram[239][3] ), .IN2(n50), .IN3(n390), .IN4(datain[3]), 
        .Q(n2159) );
  AO22X1 U167 ( .IN1(\ram[239][4] ), .IN2(n50), .IN3(n390), .IN4(datain[4]), 
        .Q(n2160) );
  AO22X1 U168 ( .IN1(\ram[239][5] ), .IN2(n50), .IN3(n390), .IN4(datain[5]), 
        .Q(n2161) );
  AO22X1 U169 ( .IN1(\ram[239][6] ), .IN2(n50), .IN3(n390), .IN4(datain[6]), 
        .Q(n2162) );
  AO22X1 U170 ( .IN1(\ram[239][7] ), .IN2(n50), .IN3(n390), .IN4(datain[7]), 
        .Q(n2163) );
  AO22X1 U173 ( .IN1(\ram[238][0] ), .IN2(n53), .IN3(n4088), .IN4(datain[0]), 
        .Q(n2164) );
  AO22X1 U174 ( .IN1(\ram[238][1] ), .IN2(n53), .IN3(n4088), .IN4(datain[1]), 
        .Q(n2165) );
  AO22X1 U175 ( .IN1(\ram[238][2] ), .IN2(n53), .IN3(n4088), .IN4(datain[2]), 
        .Q(n2166) );
  AO22X1 U176 ( .IN1(\ram[238][3] ), .IN2(n53), .IN3(n4088), .IN4(datain[3]), 
        .Q(n2167) );
  AO22X1 U177 ( .IN1(\ram[238][4] ), .IN2(n53), .IN3(n4088), .IN4(datain[4]), 
        .Q(n2168) );
  AO22X1 U178 ( .IN1(\ram[238][5] ), .IN2(n53), .IN3(n4088), .IN4(datain[5]), 
        .Q(n2169) );
  AO22X1 U179 ( .IN1(\ram[238][6] ), .IN2(n53), .IN3(n4088), .IN4(datain[6]), 
        .Q(n2170) );
  AO22X1 U180 ( .IN1(\ram[238][7] ), .IN2(n53), .IN3(n4088), .IN4(datain[7]), 
        .Q(n2171) );
  AO22X1 U183 ( .IN1(\ram[237][0] ), .IN2(n56), .IN3(n447), .IN4(datain[0]), 
        .Q(n2172) );
  AO22X1 U184 ( .IN1(\ram[237][1] ), .IN2(n56), .IN3(n447), .IN4(datain[1]), 
        .Q(n2173) );
  AO22X1 U185 ( .IN1(\ram[237][2] ), .IN2(n56), .IN3(n447), .IN4(datain[2]), 
        .Q(n2174) );
  AO22X1 U186 ( .IN1(\ram[237][3] ), .IN2(n56), .IN3(n447), .IN4(datain[3]), 
        .Q(n2175) );
  AO22X1 U187 ( .IN1(\ram[237][4] ), .IN2(n56), .IN3(n447), .IN4(datain[4]), 
        .Q(n2176) );
  AO22X1 U188 ( .IN1(\ram[237][5] ), .IN2(n56), .IN3(n447), .IN4(datain[5]), 
        .Q(n2177) );
  AO22X1 U189 ( .IN1(\ram[237][6] ), .IN2(n56), .IN3(n447), .IN4(datain[6]), 
        .Q(n2178) );
  AO22X1 U190 ( .IN1(\ram[237][7] ), .IN2(n56), .IN3(n447), .IN4(datain[7]), 
        .Q(n2179) );
  AO22X1 U193 ( .IN1(\ram[236][0] ), .IN2(n59), .IN3(n765), .IN4(datain[0]), 
        .Q(n2180) );
  AO22X1 U194 ( .IN1(\ram[236][1] ), .IN2(n59), .IN3(n765), .IN4(datain[1]), 
        .Q(n2181) );
  AO22X1 U195 ( .IN1(\ram[236][2] ), .IN2(n59), .IN3(n765), .IN4(datain[2]), 
        .Q(n2182) );
  AO22X1 U196 ( .IN1(\ram[236][3] ), .IN2(n59), .IN3(n765), .IN4(datain[3]), 
        .Q(n2183) );
  AO22X1 U197 ( .IN1(\ram[236][4] ), .IN2(n59), .IN3(n765), .IN4(datain[4]), 
        .Q(n2184) );
  AO22X1 U198 ( .IN1(\ram[236][5] ), .IN2(n59), .IN3(n765), .IN4(datain[5]), 
        .Q(n2185) );
  AO22X1 U199 ( .IN1(\ram[236][6] ), .IN2(n59), .IN3(n765), .IN4(datain[6]), 
        .Q(n2186) );
  AO22X1 U200 ( .IN1(\ram[236][7] ), .IN2(n59), .IN3(n765), .IN4(datain[7]), 
        .Q(n2187) );
  AO22X1 U203 ( .IN1(\ram[235][0] ), .IN2(n62), .IN3(n330), .IN4(datain[0]), 
        .Q(n2188) );
  AO22X1 U204 ( .IN1(\ram[235][1] ), .IN2(n62), .IN3(n330), .IN4(datain[1]), 
        .Q(n2189) );
  AO22X1 U205 ( .IN1(\ram[235][2] ), .IN2(n62), .IN3(n330), .IN4(datain[2]), 
        .Q(n2190) );
  AO22X1 U206 ( .IN1(\ram[235][3] ), .IN2(n62), .IN3(n330), .IN4(datain[3]), 
        .Q(n2191) );
  AO22X1 U207 ( .IN1(\ram[235][4] ), .IN2(n62), .IN3(n330), .IN4(datain[4]), 
        .Q(n2192) );
  AO22X1 U208 ( .IN1(\ram[235][5] ), .IN2(n62), .IN3(n330), .IN4(datain[5]), 
        .Q(n2193) );
  AO22X1 U209 ( .IN1(\ram[235][6] ), .IN2(n62), .IN3(n330), .IN4(datain[6]), 
        .Q(n2194) );
  AO22X1 U210 ( .IN1(\ram[235][7] ), .IN2(n62), .IN3(n330), .IN4(datain[7]), 
        .Q(n2195) );
  AO22X1 U213 ( .IN1(\ram[234][0] ), .IN2(n65), .IN3(n4082), .IN4(datain[0]), 
        .Q(n2196) );
  AO22X1 U214 ( .IN1(\ram[234][1] ), .IN2(n65), .IN3(n4082), .IN4(datain[1]), 
        .Q(n2197) );
  AO22X1 U215 ( .IN1(\ram[234][2] ), .IN2(n65), .IN3(n4082), .IN4(datain[2]), 
        .Q(n2198) );
  AO22X1 U216 ( .IN1(\ram[234][3] ), .IN2(n65), .IN3(n4082), .IN4(datain[3]), 
        .Q(n2199) );
  AO22X1 U217 ( .IN1(\ram[234][4] ), .IN2(n65), .IN3(n4082), .IN4(datain[4]), 
        .Q(n2200) );
  AO22X1 U218 ( .IN1(\ram[234][5] ), .IN2(n65), .IN3(n4082), .IN4(datain[5]), 
        .Q(n2201) );
  AO22X1 U219 ( .IN1(\ram[234][6] ), .IN2(n65), .IN3(n4082), .IN4(datain[6]), 
        .Q(n2202) );
  AO22X1 U220 ( .IN1(\ram[234][7] ), .IN2(n65), .IN3(n4082), .IN4(datain[7]), 
        .Q(n2203) );
  AO22X1 U223 ( .IN1(\ram[233][0] ), .IN2(n68), .IN3(n429), .IN4(datain[0]), 
        .Q(n2204) );
  AO22X1 U224 ( .IN1(\ram[233][1] ), .IN2(n68), .IN3(n429), .IN4(datain[1]), 
        .Q(n2205) );
  AO22X1 U225 ( .IN1(\ram[233][2] ), .IN2(n68), .IN3(n429), .IN4(datain[2]), 
        .Q(n2206) );
  AO22X1 U226 ( .IN1(\ram[233][3] ), .IN2(n68), .IN3(n429), .IN4(datain[3]), 
        .Q(n2207) );
  AO22X1 U227 ( .IN1(\ram[233][4] ), .IN2(n68), .IN3(n429), .IN4(datain[4]), 
        .Q(n2208) );
  AO22X1 U228 ( .IN1(\ram[233][5] ), .IN2(n68), .IN3(n429), .IN4(datain[5]), 
        .Q(n2209) );
  AO22X1 U229 ( .IN1(\ram[233][6] ), .IN2(n68), .IN3(n429), .IN4(datain[6]), 
        .Q(n2210) );
  AO22X1 U230 ( .IN1(\ram[233][7] ), .IN2(n68), .IN3(n429), .IN4(datain[7]), 
        .Q(n2211) );
  AO22X1 U233 ( .IN1(\ram[232][0] ), .IN2(n71), .IN3(n720), .IN4(datain[0]), 
        .Q(n2212) );
  AO22X1 U234 ( .IN1(\ram[232][1] ), .IN2(n71), .IN3(n720), .IN4(datain[1]), 
        .Q(n2213) );
  AO22X1 U235 ( .IN1(\ram[232][2] ), .IN2(n71), .IN3(n720), .IN4(datain[2]), 
        .Q(n2214) );
  AO22X1 U236 ( .IN1(\ram[232][3] ), .IN2(n71), .IN3(n720), .IN4(datain[3]), 
        .Q(n2215) );
  AO22X1 U237 ( .IN1(\ram[232][4] ), .IN2(n71), .IN3(n720), .IN4(datain[4]), 
        .Q(n2216) );
  AO22X1 U238 ( .IN1(\ram[232][5] ), .IN2(n71), .IN3(n720), .IN4(datain[5]), 
        .Q(n2217) );
  AO22X1 U239 ( .IN1(\ram[232][6] ), .IN2(n71), .IN3(n720), .IN4(datain[6]), 
        .Q(n2218) );
  AO22X1 U240 ( .IN1(\ram[232][7] ), .IN2(n71), .IN3(n720), .IN4(datain[7]), 
        .Q(n2219) );
  AO22X1 U243 ( .IN1(\ram[231][0] ), .IN2(n74), .IN3(n573), .IN4(datain[0]), 
        .Q(n2220) );
  AO22X1 U244 ( .IN1(\ram[231][1] ), .IN2(n74), .IN3(n573), .IN4(datain[1]), 
        .Q(n2221) );
  AO22X1 U245 ( .IN1(\ram[231][2] ), .IN2(n74), .IN3(n573), .IN4(datain[2]), 
        .Q(n2222) );
  AO22X1 U246 ( .IN1(\ram[231][3] ), .IN2(n74), .IN3(n573), .IN4(datain[3]), 
        .Q(n2223) );
  AO22X1 U247 ( .IN1(\ram[231][4] ), .IN2(n74), .IN3(n573), .IN4(datain[4]), 
        .Q(n2224) );
  AO22X1 U248 ( .IN1(\ram[231][5] ), .IN2(n74), .IN3(n573), .IN4(datain[5]), 
        .Q(n2225) );
  AO22X1 U249 ( .IN1(\ram[231][6] ), .IN2(n74), .IN3(n573), .IN4(datain[6]), 
        .Q(n2226) );
  AO22X1 U250 ( .IN1(\ram[231][7] ), .IN2(n74), .IN3(n573), .IN4(datain[7]), 
        .Q(n2227) );
  AO22X1 U253 ( .IN1(\ram[230][0] ), .IN2(n77), .IN3(n4162), .IN4(datain[0]), 
        .Q(n2228) );
  AO22X1 U254 ( .IN1(\ram[230][1] ), .IN2(n77), .IN3(n4162), .IN4(datain[1]), 
        .Q(n2229) );
  AO22X1 U255 ( .IN1(\ram[230][2] ), .IN2(n77), .IN3(n4162), .IN4(datain[2]), 
        .Q(n2230) );
  AO22X1 U256 ( .IN1(\ram[230][3] ), .IN2(n77), .IN3(n4162), .IN4(datain[3]), 
        .Q(n2231) );
  AO22X1 U257 ( .IN1(\ram[230][4] ), .IN2(n77), .IN3(n4162), .IN4(datain[4]), 
        .Q(n2232) );
  AO22X1 U258 ( .IN1(\ram[230][5] ), .IN2(n77), .IN3(n4162), .IN4(datain[5]), 
        .Q(n2233) );
  AO22X1 U259 ( .IN1(\ram[230][6] ), .IN2(n77), .IN3(n4162), .IN4(datain[6]), 
        .Q(n2234) );
  AO22X1 U260 ( .IN1(\ram[230][7] ), .IN2(n77), .IN3(n4162), .IN4(datain[7]), 
        .Q(n2235) );
  AO22X1 U263 ( .IN1(\ram[229][0] ), .IN2(n80), .IN3(n669), .IN4(datain[0]), 
        .Q(n2236) );
  AO22X1 U264 ( .IN1(\ram[229][1] ), .IN2(n80), .IN3(n669), .IN4(datain[1]), 
        .Q(n2237) );
  AO22X1 U265 ( .IN1(\ram[229][2] ), .IN2(n80), .IN3(n669), .IN4(datain[2]), 
        .Q(n2238) );
  AO22X1 U266 ( .IN1(\ram[229][3] ), .IN2(n80), .IN3(n669), .IN4(datain[3]), 
        .Q(n2239) );
  AO22X1 U267 ( .IN1(\ram[229][4] ), .IN2(n80), .IN3(n669), .IN4(datain[4]), 
        .Q(n2240) );
  AO22X1 U268 ( .IN1(\ram[229][5] ), .IN2(n80), .IN3(n669), .IN4(datain[5]), 
        .Q(n2241) );
  AO22X1 U269 ( .IN1(\ram[229][6] ), .IN2(n80), .IN3(n669), .IN4(datain[6]), 
        .Q(n2242) );
  AO22X1 U270 ( .IN1(\ram[229][7] ), .IN2(n80), .IN3(n669), .IN4(datain[7]), 
        .Q(n2243) );
  AO22X1 U273 ( .IN1(\ram[228][0] ), .IN2(n83), .IN3(n4114), .IN4(datain[0]), 
        .Q(n2244) );
  AO22X1 U274 ( .IN1(\ram[228][1] ), .IN2(n83), .IN3(n4114), .IN4(datain[1]), 
        .Q(n2245) );
  AO22X1 U275 ( .IN1(\ram[228][2] ), .IN2(n83), .IN3(n4114), .IN4(datain[2]), 
        .Q(n2246) );
  AO22X1 U276 ( .IN1(\ram[228][3] ), .IN2(n83), .IN3(n4114), .IN4(datain[3]), 
        .Q(n2247) );
  AO22X1 U277 ( .IN1(\ram[228][4] ), .IN2(n83), .IN3(n4114), .IN4(datain[4]), 
        .Q(n2248) );
  AO22X1 U278 ( .IN1(\ram[228][5] ), .IN2(n83), .IN3(n4114), .IN4(datain[5]), 
        .Q(n2249) );
  AO22X1 U279 ( .IN1(\ram[228][6] ), .IN2(n83), .IN3(n4114), .IN4(datain[6]), 
        .Q(n2250) );
  AO22X1 U280 ( .IN1(\ram[228][7] ), .IN2(n83), .IN3(n4114), .IN4(datain[7]), 
        .Q(n2251) );
  AO22X1 U283 ( .IN1(\ram[227][0] ), .IN2(n86), .IN3(n525), .IN4(datain[0]), 
        .Q(n2252) );
  AO22X1 U284 ( .IN1(\ram[227][1] ), .IN2(n86), .IN3(n525), .IN4(datain[1]), 
        .Q(n2253) );
  AO22X1 U285 ( .IN1(\ram[227][2] ), .IN2(n86), .IN3(n525), .IN4(datain[2]), 
        .Q(n2254) );
  AO22X1 U286 ( .IN1(\ram[227][3] ), .IN2(n86), .IN3(n525), .IN4(datain[3]), 
        .Q(n2255) );
  AO22X1 U287 ( .IN1(\ram[227][4] ), .IN2(n86), .IN3(n525), .IN4(datain[4]), 
        .Q(n2256) );
  AO22X1 U288 ( .IN1(\ram[227][5] ), .IN2(n86), .IN3(n525), .IN4(datain[5]), 
        .Q(n2257) );
  AO22X1 U289 ( .IN1(\ram[227][6] ), .IN2(n86), .IN3(n525), .IN4(datain[6]), 
        .Q(n2258) );
  AO22X1 U290 ( .IN1(\ram[227][7] ), .IN2(n86), .IN3(n525), .IN4(datain[7]), 
        .Q(n2259) );
  AO22X1 U293 ( .IN1(\ram[226][0] ), .IN2(n89), .IN3(n4145), .IN4(datain[0]), 
        .Q(n2260) );
  AO22X1 U294 ( .IN1(\ram[226][1] ), .IN2(n89), .IN3(n4145), .IN4(datain[1]), 
        .Q(n2261) );
  AO22X1 U295 ( .IN1(\ram[226][2] ), .IN2(n89), .IN3(n4145), .IN4(datain[2]), 
        .Q(n2262) );
  AO22X1 U296 ( .IN1(\ram[226][3] ), .IN2(n89), .IN3(n4145), .IN4(datain[3]), 
        .Q(n2263) );
  AO22X1 U297 ( .IN1(\ram[226][4] ), .IN2(n89), .IN3(n4145), .IN4(datain[4]), 
        .Q(n2264) );
  AO22X1 U298 ( .IN1(\ram[226][5] ), .IN2(n89), .IN3(n4145), .IN4(datain[5]), 
        .Q(n2265) );
  AO22X1 U299 ( .IN1(\ram[226][6] ), .IN2(n89), .IN3(n4145), .IN4(datain[6]), 
        .Q(n2266) );
  AO22X1 U300 ( .IN1(\ram[226][7] ), .IN2(n89), .IN3(n4145), .IN4(datain[7]), 
        .Q(n2267) );
  AO22X1 U303 ( .IN1(\ram[225][0] ), .IN2(n92), .IN3(n621), .IN4(datain[0]), 
        .Q(n2268) );
  AO22X1 U304 ( .IN1(\ram[225][1] ), .IN2(n92), .IN3(n621), .IN4(datain[1]), 
        .Q(n2269) );
  AO22X1 U305 ( .IN1(\ram[225][2] ), .IN2(n92), .IN3(n621), .IN4(datain[2]), 
        .Q(n2270) );
  AO22X1 U306 ( .IN1(\ram[225][3] ), .IN2(n92), .IN3(n621), .IN4(datain[3]), 
        .Q(n2271) );
  AO22X1 U307 ( .IN1(\ram[225][4] ), .IN2(n92), .IN3(n621), .IN4(datain[4]), 
        .Q(n2272) );
  AO22X1 U308 ( .IN1(\ram[225][5] ), .IN2(n92), .IN3(n621), .IN4(datain[5]), 
        .Q(n2273) );
  AO22X1 U309 ( .IN1(\ram[225][6] ), .IN2(n92), .IN3(n621), .IN4(datain[6]), 
        .Q(n2274) );
  AO22X1 U310 ( .IN1(\ram[225][7] ), .IN2(n92), .IN3(n621), .IN4(datain[7]), 
        .Q(n2275) );
  AO22X1 U313 ( .IN1(\ram[224][0] ), .IN2(n95), .IN3(n4127), .IN4(datain[0]), 
        .Q(n2276) );
  AO22X1 U314 ( .IN1(\ram[224][1] ), .IN2(n95), .IN3(n4127), .IN4(datain[1]), 
        .Q(n2277) );
  AO22X1 U315 ( .IN1(\ram[224][2] ), .IN2(n95), .IN3(n4127), .IN4(datain[2]), 
        .Q(n2278) );
  AO22X1 U316 ( .IN1(\ram[224][3] ), .IN2(n95), .IN3(n4127), .IN4(datain[3]), 
        .Q(n2279) );
  AO22X1 U317 ( .IN1(\ram[224][4] ), .IN2(n95), .IN3(n4127), .IN4(datain[4]), 
        .Q(n2280) );
  AO22X1 U318 ( .IN1(\ram[224][5] ), .IN2(n95), .IN3(n4127), .IN4(datain[5]), 
        .Q(n2281) );
  AO22X1 U319 ( .IN1(\ram[224][6] ), .IN2(n95), .IN3(n4127), .IN4(datain[6]), 
        .Q(n2282) );
  AO22X1 U320 ( .IN1(\ram[224][7] ), .IN2(n95), .IN3(n4127), .IN4(datain[7]), 
        .Q(n2283) );
  AO22X1 U323 ( .IN1(\ram[223][0] ), .IN2(n98), .IN3(n372), .IN4(datain[0]), 
        .Q(n2284) );
  AO22X1 U324 ( .IN1(\ram[223][1] ), .IN2(n98), .IN3(n372), .IN4(datain[1]), 
        .Q(n2285) );
  AO22X1 U325 ( .IN1(\ram[223][2] ), .IN2(n98), .IN3(n372), .IN4(datain[2]), 
        .Q(n2286) );
  AO22X1 U326 ( .IN1(\ram[223][3] ), .IN2(n98), .IN3(n372), .IN4(datain[3]), 
        .Q(n2287) );
  AO22X1 U327 ( .IN1(\ram[223][4] ), .IN2(n98), .IN3(n372), .IN4(datain[4]), 
        .Q(n2288) );
  AO22X1 U328 ( .IN1(\ram[223][5] ), .IN2(n98), .IN3(n372), .IN4(datain[5]), 
        .Q(n2289) );
  AO22X1 U329 ( .IN1(\ram[223][6] ), .IN2(n98), .IN3(n372), .IN4(datain[6]), 
        .Q(n2290) );
  AO22X1 U330 ( .IN1(\ram[223][7] ), .IN2(n98), .IN3(n372), .IN4(datain[7]), 
        .Q(n2291) );
  AO22X1 U333 ( .IN1(\ram[222][0] ), .IN2(n101), .IN3(n4098), .IN4(datain[0]), 
        .Q(n2292) );
  AO22X1 U334 ( .IN1(\ram[222][1] ), .IN2(n101), .IN3(n4098), .IN4(datain[1]), 
        .Q(n2293) );
  AO22X1 U335 ( .IN1(\ram[222][2] ), .IN2(n101), .IN3(n4098), .IN4(datain[2]), 
        .Q(n2294) );
  AO22X1 U336 ( .IN1(\ram[222][3] ), .IN2(n101), .IN3(n4098), .IN4(datain[3]), 
        .Q(n2295) );
  AO22X1 U337 ( .IN1(\ram[222][4] ), .IN2(n101), .IN3(n4098), .IN4(datain[4]), 
        .Q(n2296) );
  AO22X1 U338 ( .IN1(\ram[222][5] ), .IN2(n101), .IN3(n4098), .IN4(datain[5]), 
        .Q(n2297) );
  AO22X1 U339 ( .IN1(\ram[222][6] ), .IN2(n101), .IN3(n4098), .IN4(datain[6]), 
        .Q(n2298) );
  AO22X1 U340 ( .IN1(\ram[222][7] ), .IN2(n101), .IN3(n4098), .IN4(datain[7]), 
        .Q(n2299) );
  AO22X1 U343 ( .IN1(\ram[221][0] ), .IN2(n104), .IN3(n477), .IN4(datain[0]), 
        .Q(n2300) );
  AO22X1 U344 ( .IN1(\ram[221][1] ), .IN2(n104), .IN3(n477), .IN4(datain[1]), 
        .Q(n2301) );
  AO22X1 U345 ( .IN1(\ram[221][2] ), .IN2(n104), .IN3(n477), .IN4(datain[2]), 
        .Q(n2302) );
  AO22X1 U346 ( .IN1(\ram[221][3] ), .IN2(n104), .IN3(n477), .IN4(datain[3]), 
        .Q(n2303) );
  AO22X1 U347 ( .IN1(\ram[221][4] ), .IN2(n104), .IN3(n477), .IN4(datain[4]), 
        .Q(n2304) );
  AO22X1 U348 ( .IN1(\ram[221][5] ), .IN2(n104), .IN3(n477), .IN4(datain[5]), 
        .Q(n2305) );
  AO22X1 U349 ( .IN1(\ram[221][6] ), .IN2(n104), .IN3(n477), .IN4(datain[6]), 
        .Q(n2306) );
  AO22X1 U350 ( .IN1(\ram[221][7] ), .IN2(n104), .IN3(n477), .IN4(datain[7]), 
        .Q(n2307) );
  AO22X1 U353 ( .IN1(\ram[220][0] ), .IN2(n107), .IN3(n759), .IN4(datain[0]), 
        .Q(n2308) );
  AO22X1 U354 ( .IN1(\ram[220][1] ), .IN2(n107), .IN3(n759), .IN4(datain[1]), 
        .Q(n2309) );
  AO22X1 U355 ( .IN1(\ram[220][2] ), .IN2(n107), .IN3(n759), .IN4(datain[2]), 
        .Q(n2310) );
  AO22X1 U356 ( .IN1(\ram[220][3] ), .IN2(n107), .IN3(n759), .IN4(datain[3]), 
        .Q(n2311) );
  AO22X1 U357 ( .IN1(\ram[220][4] ), .IN2(n107), .IN3(n759), .IN4(datain[4]), 
        .Q(n2312) );
  AO22X1 U358 ( .IN1(\ram[220][5] ), .IN2(n107), .IN3(n759), .IN4(datain[5]), 
        .Q(n2313) );
  AO22X1 U359 ( .IN1(\ram[220][6] ), .IN2(n107), .IN3(n759), .IN4(datain[6]), 
        .Q(n2314) );
  AO22X1 U360 ( .IN1(\ram[220][7] ), .IN2(n107), .IN3(n759), .IN4(datain[7]), 
        .Q(n2315) );
  AO22X1 U363 ( .IN1(\ram[219][0] ), .IN2(n110), .IN3(n324), .IN4(datain[0]), 
        .Q(n2316) );
  AO22X1 U364 ( .IN1(\ram[219][1] ), .IN2(n110), .IN3(n324), .IN4(datain[1]), 
        .Q(n2317) );
  AO22X1 U365 ( .IN1(\ram[219][2] ), .IN2(n110), .IN3(n324), .IN4(datain[2]), 
        .Q(n2318) );
  AO22X1 U366 ( .IN1(\ram[219][3] ), .IN2(n110), .IN3(n324), .IN4(datain[3]), 
        .Q(n2319) );
  AO22X1 U367 ( .IN1(\ram[219][4] ), .IN2(n110), .IN3(n324), .IN4(datain[4]), 
        .Q(n2320) );
  AO22X1 U368 ( .IN1(\ram[219][5] ), .IN2(n110), .IN3(n324), .IN4(datain[5]), 
        .Q(n2321) );
  AO22X1 U369 ( .IN1(\ram[219][6] ), .IN2(n110), .IN3(n324), .IN4(datain[6]), 
        .Q(n2322) );
  AO22X1 U370 ( .IN1(\ram[219][7] ), .IN2(n110), .IN3(n324), .IN4(datain[7]), 
        .Q(n2323) );
  AO22X1 U373 ( .IN1(\ram[218][0] ), .IN2(n113), .IN3(n4080), .IN4(datain[0]), 
        .Q(n2324) );
  AO22X1 U374 ( .IN1(\ram[218][1] ), .IN2(n113), .IN3(n4080), .IN4(datain[1]), 
        .Q(n2325) );
  AO22X1 U375 ( .IN1(\ram[218][2] ), .IN2(n113), .IN3(n4080), .IN4(datain[2]), 
        .Q(n2326) );
  AO22X1 U376 ( .IN1(\ram[218][3] ), .IN2(n113), .IN3(n4080), .IN4(datain[3]), 
        .Q(n2327) );
  AO22X1 U377 ( .IN1(\ram[218][4] ), .IN2(n113), .IN3(n4080), .IN4(datain[4]), 
        .Q(n2328) );
  AO22X1 U378 ( .IN1(\ram[218][5] ), .IN2(n113), .IN3(n4080), .IN4(datain[5]), 
        .Q(n2329) );
  AO22X1 U379 ( .IN1(\ram[218][6] ), .IN2(n113), .IN3(n4080), .IN4(datain[6]), 
        .Q(n2330) );
  AO22X1 U380 ( .IN1(\ram[218][7] ), .IN2(n113), .IN3(n4080), .IN4(datain[7]), 
        .Q(n2331) );
  AO22X1 U383 ( .IN1(\ram[217][0] ), .IN2(n116), .IN3(n423), .IN4(datain[0]), 
        .Q(n2332) );
  AO22X1 U384 ( .IN1(\ram[217][1] ), .IN2(n116), .IN3(n423), .IN4(datain[1]), 
        .Q(n2333) );
  AO22X1 U385 ( .IN1(\ram[217][2] ), .IN2(n116), .IN3(n423), .IN4(datain[2]), 
        .Q(n2334) );
  AO22X1 U386 ( .IN1(\ram[217][3] ), .IN2(n116), .IN3(n423), .IN4(datain[3]), 
        .Q(n2335) );
  AO22X1 U387 ( .IN1(\ram[217][4] ), .IN2(n116), .IN3(n423), .IN4(datain[4]), 
        .Q(n2336) );
  AO22X1 U388 ( .IN1(\ram[217][5] ), .IN2(n116), .IN3(n423), .IN4(datain[5]), 
        .Q(n2337) );
  AO22X1 U389 ( .IN1(\ram[217][6] ), .IN2(n116), .IN3(n423), .IN4(datain[6]), 
        .Q(n2338) );
  AO22X1 U390 ( .IN1(\ram[217][7] ), .IN2(n116), .IN3(n423), .IN4(datain[7]), 
        .Q(n2339) );
  AO22X1 U393 ( .IN1(\ram[216][0] ), .IN2(n119), .IN3(n711), .IN4(datain[0]), 
        .Q(n2340) );
  AO22X1 U394 ( .IN1(\ram[216][1] ), .IN2(n119), .IN3(n711), .IN4(datain[1]), 
        .Q(n2341) );
  AO22X1 U395 ( .IN1(\ram[216][2] ), .IN2(n119), .IN3(n711), .IN4(datain[2]), 
        .Q(n2342) );
  AO22X1 U396 ( .IN1(\ram[216][3] ), .IN2(n119), .IN3(n711), .IN4(datain[3]), 
        .Q(n2343) );
  AO22X1 U397 ( .IN1(\ram[216][4] ), .IN2(n119), .IN3(n711), .IN4(datain[4]), 
        .Q(n2344) );
  AO22X1 U398 ( .IN1(\ram[216][5] ), .IN2(n119), .IN3(n711), .IN4(datain[5]), 
        .Q(n2345) );
  AO22X1 U399 ( .IN1(\ram[216][6] ), .IN2(n119), .IN3(n711), .IN4(datain[6]), 
        .Q(n2346) );
  AO22X1 U400 ( .IN1(\ram[216][7] ), .IN2(n119), .IN3(n711), .IN4(datain[7]), 
        .Q(n2347) );
  AO22X1 U403 ( .IN1(\ram[215][0] ), .IN2(n122), .IN3(n564), .IN4(datain[0]), 
        .Q(n2348) );
  AO22X1 U404 ( .IN1(\ram[215][1] ), .IN2(n122), .IN3(n564), .IN4(datain[1]), 
        .Q(n2349) );
  AO22X1 U405 ( .IN1(\ram[215][2] ), .IN2(n122), .IN3(n564), .IN4(datain[2]), 
        .Q(n2350) );
  AO22X1 U406 ( .IN1(\ram[215][3] ), .IN2(n122), .IN3(n564), .IN4(datain[3]), 
        .Q(n2351) );
  AO22X1 U407 ( .IN1(\ram[215][4] ), .IN2(n122), .IN3(n564), .IN4(datain[4]), 
        .Q(n2352) );
  AO22X1 U408 ( .IN1(\ram[215][5] ), .IN2(n122), .IN3(n564), .IN4(datain[5]), 
        .Q(n2353) );
  AO22X1 U409 ( .IN1(\ram[215][6] ), .IN2(n122), .IN3(n564), .IN4(datain[6]), 
        .Q(n2354) );
  AO22X1 U410 ( .IN1(\ram[215][7] ), .IN2(n122), .IN3(n564), .IN4(datain[7]), 
        .Q(n2355) );
  AO22X1 U413 ( .IN1(\ram[214][0] ), .IN2(n125), .IN3(n4159), .IN4(datain[0]), 
        .Q(n2356) );
  AO22X1 U414 ( .IN1(\ram[214][1] ), .IN2(n125), .IN3(n4159), .IN4(datain[1]), 
        .Q(n2357) );
  AO22X1 U415 ( .IN1(\ram[214][2] ), .IN2(n125), .IN3(n4159), .IN4(datain[2]), 
        .Q(n2358) );
  AO22X1 U416 ( .IN1(\ram[214][3] ), .IN2(n125), .IN3(n4159), .IN4(datain[3]), 
        .Q(n2359) );
  AO22X1 U417 ( .IN1(\ram[214][4] ), .IN2(n125), .IN3(n4159), .IN4(datain[4]), 
        .Q(n2360) );
  AO22X1 U418 ( .IN1(\ram[214][5] ), .IN2(n125), .IN3(n4159), .IN4(datain[5]), 
        .Q(n2361) );
  AO22X1 U419 ( .IN1(\ram[214][6] ), .IN2(n125), .IN3(n4159), .IN4(datain[6]), 
        .Q(n2362) );
  AO22X1 U420 ( .IN1(\ram[214][7] ), .IN2(n125), .IN3(n4159), .IN4(datain[7]), 
        .Q(n2363) );
  AO22X1 U423 ( .IN1(\ram[213][0] ), .IN2(n128), .IN3(n660), .IN4(datain[0]), 
        .Q(n2364) );
  AO22X1 U424 ( .IN1(\ram[213][1] ), .IN2(n128), .IN3(n660), .IN4(datain[1]), 
        .Q(n2365) );
  AO22X1 U425 ( .IN1(\ram[213][2] ), .IN2(n128), .IN3(n660), .IN4(datain[2]), 
        .Q(n2366) );
  AO22X1 U426 ( .IN1(\ram[213][3] ), .IN2(n128), .IN3(n660), .IN4(datain[3]), 
        .Q(n2367) );
  AO22X1 U427 ( .IN1(\ram[213][4] ), .IN2(n128), .IN3(n660), .IN4(datain[4]), 
        .Q(n2368) );
  AO22X1 U428 ( .IN1(\ram[213][5] ), .IN2(n128), .IN3(n660), .IN4(datain[5]), 
        .Q(n2369) );
  AO22X1 U429 ( .IN1(\ram[213][6] ), .IN2(n128), .IN3(n660), .IN4(datain[6]), 
        .Q(n2370) );
  AO22X1 U430 ( .IN1(\ram[213][7] ), .IN2(n128), .IN3(n660), .IN4(datain[7]), 
        .Q(n2371) );
  AO22X1 U433 ( .IN1(\ram[212][0] ), .IN2(n131), .IN3(n4111), .IN4(datain[0]), 
        .Q(n2372) );
  AO22X1 U434 ( .IN1(\ram[212][1] ), .IN2(n131), .IN3(n4111), .IN4(datain[1]), 
        .Q(n2373) );
  AO22X1 U435 ( .IN1(\ram[212][2] ), .IN2(n131), .IN3(n4111), .IN4(datain[2]), 
        .Q(n2374) );
  AO22X1 U436 ( .IN1(\ram[212][3] ), .IN2(n131), .IN3(n4111), .IN4(datain[3]), 
        .Q(n2375) );
  AO22X1 U437 ( .IN1(\ram[212][4] ), .IN2(n131), .IN3(n4111), .IN4(datain[4]), 
        .Q(n2376) );
  AO22X1 U438 ( .IN1(\ram[212][5] ), .IN2(n131), .IN3(n4111), .IN4(datain[5]), 
        .Q(n2377) );
  AO22X1 U439 ( .IN1(\ram[212][6] ), .IN2(n131), .IN3(n4111), .IN4(datain[6]), 
        .Q(n2378) );
  AO22X1 U440 ( .IN1(\ram[212][7] ), .IN2(n131), .IN3(n4111), .IN4(datain[7]), 
        .Q(n2379) );
  AO22X1 U443 ( .IN1(\ram[211][0] ), .IN2(n134), .IN3(n516), .IN4(datain[0]), 
        .Q(n2380) );
  AO22X1 U444 ( .IN1(\ram[211][1] ), .IN2(n134), .IN3(n516), .IN4(datain[1]), 
        .Q(n2381) );
  AO22X1 U445 ( .IN1(\ram[211][2] ), .IN2(n134), .IN3(n516), .IN4(datain[2]), 
        .Q(n2382) );
  AO22X1 U446 ( .IN1(\ram[211][3] ), .IN2(n134), .IN3(n516), .IN4(datain[3]), 
        .Q(n2383) );
  AO22X1 U447 ( .IN1(\ram[211][4] ), .IN2(n134), .IN3(n516), .IN4(datain[4]), 
        .Q(n2384) );
  AO22X1 U448 ( .IN1(\ram[211][5] ), .IN2(n134), .IN3(n516), .IN4(datain[5]), 
        .Q(n2385) );
  AO22X1 U449 ( .IN1(\ram[211][6] ), .IN2(n134), .IN3(n516), .IN4(datain[6]), 
        .Q(n2386) );
  AO22X1 U450 ( .IN1(\ram[211][7] ), .IN2(n134), .IN3(n516), .IN4(datain[7]), 
        .Q(n2387) );
  AO22X1 U453 ( .IN1(\ram[210][0] ), .IN2(n137), .IN3(n4146), .IN4(datain[0]), 
        .Q(n2388) );
  AO22X1 U454 ( .IN1(\ram[210][1] ), .IN2(n137), .IN3(n4146), .IN4(datain[1]), 
        .Q(n2389) );
  AO22X1 U455 ( .IN1(\ram[210][2] ), .IN2(n137), .IN3(n4146), .IN4(datain[2]), 
        .Q(n2390) );
  AO22X1 U456 ( .IN1(\ram[210][3] ), .IN2(n137), .IN3(n4146), .IN4(datain[3]), 
        .Q(n2391) );
  AO22X1 U457 ( .IN1(\ram[210][4] ), .IN2(n137), .IN3(n4146), .IN4(datain[4]), 
        .Q(n2392) );
  AO22X1 U458 ( .IN1(\ram[210][5] ), .IN2(n137), .IN3(n4146), .IN4(datain[5]), 
        .Q(n2393) );
  AO22X1 U459 ( .IN1(\ram[210][6] ), .IN2(n137), .IN3(n4146), .IN4(datain[6]), 
        .Q(n2394) );
  AO22X1 U460 ( .IN1(\ram[210][7] ), .IN2(n137), .IN3(n4146), .IN4(datain[7]), 
        .Q(n2395) );
  AO22X1 U463 ( .IN1(\ram[209][0] ), .IN2(n140), .IN3(n612), .IN4(datain[0]), 
        .Q(n2396) );
  AO22X1 U464 ( .IN1(\ram[209][1] ), .IN2(n140), .IN3(n612), .IN4(datain[1]), 
        .Q(n2397) );
  AO22X1 U465 ( .IN1(\ram[209][2] ), .IN2(n140), .IN3(n612), .IN4(datain[2]), 
        .Q(n2398) );
  AO22X1 U466 ( .IN1(\ram[209][3] ), .IN2(n140), .IN3(n612), .IN4(datain[3]), 
        .Q(n2399) );
  AO22X1 U467 ( .IN1(\ram[209][4] ), .IN2(n140), .IN3(n612), .IN4(datain[4]), 
        .Q(n2400) );
  AO22X1 U468 ( .IN1(\ram[209][5] ), .IN2(n140), .IN3(n612), .IN4(datain[5]), 
        .Q(n2401) );
  AO22X1 U469 ( .IN1(\ram[209][6] ), .IN2(n140), .IN3(n612), .IN4(datain[6]), 
        .Q(n2402) );
  AO22X1 U470 ( .IN1(\ram[209][7] ), .IN2(n140), .IN3(n612), .IN4(datain[7]), 
        .Q(n2403) );
  AO22X1 U473 ( .IN1(\ram[208][0] ), .IN2(n143), .IN3(n4128), .IN4(datain[0]), 
        .Q(n2404) );
  AO22X1 U474 ( .IN1(\ram[208][1] ), .IN2(n143), .IN3(n4128), .IN4(datain[1]), 
        .Q(n2405) );
  AO22X1 U475 ( .IN1(\ram[208][2] ), .IN2(n143), .IN3(n4128), .IN4(datain[2]), 
        .Q(n2406) );
  AO22X1 U476 ( .IN1(\ram[208][3] ), .IN2(n143), .IN3(n4128), .IN4(datain[3]), 
        .Q(n2407) );
  AO22X1 U477 ( .IN1(\ram[208][4] ), .IN2(n143), .IN3(n4128), .IN4(datain[4]), 
        .Q(n2408) );
  AO22X1 U478 ( .IN1(\ram[208][5] ), .IN2(n143), .IN3(n4128), .IN4(datain[5]), 
        .Q(n2409) );
  AO22X1 U479 ( .IN1(\ram[208][6] ), .IN2(n143), .IN3(n4128), .IN4(datain[6]), 
        .Q(n2410) );
  AO22X1 U480 ( .IN1(\ram[208][7] ), .IN2(n143), .IN3(n4128), .IN4(datain[7]), 
        .Q(n2411) );
  AO22X1 U483 ( .IN1(\ram[207][0] ), .IN2(n146), .IN3(n375), .IN4(datain[0]), 
        .Q(n2412) );
  AO22X1 U484 ( .IN1(\ram[207][1] ), .IN2(n146), .IN3(n375), .IN4(datain[1]), 
        .Q(n2413) );
  AO22X1 U485 ( .IN1(\ram[207][2] ), .IN2(n146), .IN3(n375), .IN4(datain[2]), 
        .Q(n2414) );
  AO22X1 U486 ( .IN1(\ram[207][3] ), .IN2(n146), .IN3(n375), .IN4(datain[3]), 
        .Q(n2415) );
  AO22X1 U487 ( .IN1(\ram[207][4] ), .IN2(n146), .IN3(n375), .IN4(datain[4]), 
        .Q(n2416) );
  AO22X1 U488 ( .IN1(\ram[207][5] ), .IN2(n146), .IN3(n375), .IN4(datain[5]), 
        .Q(n2417) );
  AO22X1 U489 ( .IN1(\ram[207][6] ), .IN2(n146), .IN3(n375), .IN4(datain[6]), 
        .Q(n2418) );
  AO22X1 U490 ( .IN1(\ram[207][7] ), .IN2(n146), .IN3(n375), .IN4(datain[7]), 
        .Q(n2419) );
  AO22X1 U493 ( .IN1(\ram[206][0] ), .IN2(n149), .IN3(n4099), .IN4(datain[0]), 
        .Q(n2420) );
  AO22X1 U494 ( .IN1(\ram[206][1] ), .IN2(n149), .IN3(n4099), .IN4(datain[1]), 
        .Q(n2421) );
  AO22X1 U495 ( .IN1(\ram[206][2] ), .IN2(n149), .IN3(n4099), .IN4(datain[2]), 
        .Q(n2422) );
  AO22X1 U496 ( .IN1(\ram[206][3] ), .IN2(n149), .IN3(n4099), .IN4(datain[3]), 
        .Q(n2423) );
  AO22X1 U497 ( .IN1(\ram[206][4] ), .IN2(n149), .IN3(n4099), .IN4(datain[4]), 
        .Q(n2424) );
  AO22X1 U498 ( .IN1(\ram[206][5] ), .IN2(n149), .IN3(n4099), .IN4(datain[5]), 
        .Q(n2425) );
  AO22X1 U499 ( .IN1(\ram[206][6] ), .IN2(n149), .IN3(n4099), .IN4(datain[6]), 
        .Q(n2426) );
  AO22X1 U500 ( .IN1(\ram[206][7] ), .IN2(n149), .IN3(n4099), .IN4(datain[7]), 
        .Q(n2427) );
  AO22X1 U503 ( .IN1(\ram[205][0] ), .IN2(n152), .IN3(n480), .IN4(datain[0]), 
        .Q(n2428) );
  AO22X1 U504 ( .IN1(\ram[205][1] ), .IN2(n152), .IN3(n480), .IN4(datain[1]), 
        .Q(n2429) );
  AO22X1 U505 ( .IN1(\ram[205][2] ), .IN2(n152), .IN3(n480), .IN4(datain[2]), 
        .Q(n2430) );
  AO22X1 U506 ( .IN1(\ram[205][3] ), .IN2(n152), .IN3(n480), .IN4(datain[3]), 
        .Q(n2431) );
  AO22X1 U507 ( .IN1(\ram[205][4] ), .IN2(n152), .IN3(n480), .IN4(datain[4]), 
        .Q(n2432) );
  AO22X1 U508 ( .IN1(\ram[205][5] ), .IN2(n152), .IN3(n480), .IN4(datain[5]), 
        .Q(n2433) );
  AO22X1 U509 ( .IN1(\ram[205][6] ), .IN2(n152), .IN3(n480), .IN4(datain[6]), 
        .Q(n2434) );
  AO22X1 U510 ( .IN1(\ram[205][7] ), .IN2(n152), .IN3(n480), .IN4(datain[7]), 
        .Q(n2435) );
  AO22X1 U513 ( .IN1(\ram[204][0] ), .IN2(n155), .IN3(n762), .IN4(datain[0]), 
        .Q(n2436) );
  AO22X1 U514 ( .IN1(\ram[204][1] ), .IN2(n155), .IN3(n762), .IN4(datain[1]), 
        .Q(n2437) );
  AO22X1 U515 ( .IN1(\ram[204][2] ), .IN2(n155), .IN3(n762), .IN4(datain[2]), 
        .Q(n2438) );
  AO22X1 U516 ( .IN1(\ram[204][3] ), .IN2(n155), .IN3(n762), .IN4(datain[3]), 
        .Q(n2439) );
  AO22X1 U517 ( .IN1(\ram[204][4] ), .IN2(n155), .IN3(n762), .IN4(datain[4]), 
        .Q(n2440) );
  AO22X1 U518 ( .IN1(\ram[204][5] ), .IN2(n155), .IN3(n762), .IN4(datain[5]), 
        .Q(n2441) );
  AO22X1 U519 ( .IN1(\ram[204][6] ), .IN2(n155), .IN3(n762), .IN4(datain[6]), 
        .Q(n2442) );
  AO22X1 U520 ( .IN1(\ram[204][7] ), .IN2(n155), .IN3(n762), .IN4(datain[7]), 
        .Q(n2443) );
  AO22X1 U523 ( .IN1(\ram[203][0] ), .IN2(n158), .IN3(n327), .IN4(datain[0]), 
        .Q(n2444) );
  AO22X1 U524 ( .IN1(\ram[203][1] ), .IN2(n158), .IN3(n327), .IN4(datain[1]), 
        .Q(n2445) );
  AO22X1 U525 ( .IN1(\ram[203][2] ), .IN2(n158), .IN3(n327), .IN4(datain[2]), 
        .Q(n2446) );
  AO22X1 U526 ( .IN1(\ram[203][3] ), .IN2(n158), .IN3(n327), .IN4(datain[3]), 
        .Q(n2447) );
  AO22X1 U527 ( .IN1(\ram[203][4] ), .IN2(n158), .IN3(n327), .IN4(datain[4]), 
        .Q(n2448) );
  AO22X1 U528 ( .IN1(\ram[203][5] ), .IN2(n158), .IN3(n327), .IN4(datain[5]), 
        .Q(n2449) );
  AO22X1 U529 ( .IN1(\ram[203][6] ), .IN2(n158), .IN3(n327), .IN4(datain[6]), 
        .Q(n2450) );
  AO22X1 U530 ( .IN1(\ram[203][7] ), .IN2(n158), .IN3(n327), .IN4(datain[7]), 
        .Q(n2451) );
  AO22X1 U533 ( .IN1(\ram[202][0] ), .IN2(n161), .IN3(n4081), .IN4(datain[0]), 
        .Q(n2452) );
  AO22X1 U534 ( .IN1(\ram[202][1] ), .IN2(n161), .IN3(n4081), .IN4(datain[1]), 
        .Q(n2453) );
  AO22X1 U535 ( .IN1(\ram[202][2] ), .IN2(n161), .IN3(n4081), .IN4(datain[2]), 
        .Q(n2454) );
  AO22X1 U536 ( .IN1(\ram[202][3] ), .IN2(n161), .IN3(n4081), .IN4(datain[3]), 
        .Q(n2455) );
  AO22X1 U537 ( .IN1(\ram[202][4] ), .IN2(n161), .IN3(n4081), .IN4(datain[4]), 
        .Q(n2456) );
  AO22X1 U538 ( .IN1(\ram[202][5] ), .IN2(n161), .IN3(n4081), .IN4(datain[5]), 
        .Q(n2457) );
  AO22X1 U539 ( .IN1(\ram[202][6] ), .IN2(n161), .IN3(n4081), .IN4(datain[6]), 
        .Q(n2458) );
  AO22X1 U540 ( .IN1(\ram[202][7] ), .IN2(n161), .IN3(n4081), .IN4(datain[7]), 
        .Q(n2459) );
  AO22X1 U543 ( .IN1(\ram[201][0] ), .IN2(n164), .IN3(n426), .IN4(datain[0]), 
        .Q(n2460) );
  AO22X1 U544 ( .IN1(\ram[201][1] ), .IN2(n164), .IN3(n426), .IN4(datain[1]), 
        .Q(n2461) );
  AO22X1 U545 ( .IN1(\ram[201][2] ), .IN2(n164), .IN3(n426), .IN4(datain[2]), 
        .Q(n2462) );
  AO22X1 U546 ( .IN1(\ram[201][3] ), .IN2(n164), .IN3(n426), .IN4(datain[3]), 
        .Q(n2463) );
  AO22X1 U547 ( .IN1(\ram[201][4] ), .IN2(n164), .IN3(n426), .IN4(datain[4]), 
        .Q(n2464) );
  AO22X1 U548 ( .IN1(\ram[201][5] ), .IN2(n164), .IN3(n426), .IN4(datain[5]), 
        .Q(n2465) );
  AO22X1 U549 ( .IN1(\ram[201][6] ), .IN2(n164), .IN3(n426), .IN4(datain[6]), 
        .Q(n2466) );
  AO22X1 U550 ( .IN1(\ram[201][7] ), .IN2(n164), .IN3(n426), .IN4(datain[7]), 
        .Q(n2467) );
  AO22X1 U553 ( .IN1(\ram[200][0] ), .IN2(n167), .IN3(n714), .IN4(datain[0]), 
        .Q(n2468) );
  AO22X1 U554 ( .IN1(\ram[200][1] ), .IN2(n167), .IN3(n714), .IN4(datain[1]), 
        .Q(n2469) );
  AO22X1 U555 ( .IN1(\ram[200][2] ), .IN2(n167), .IN3(n714), .IN4(datain[2]), 
        .Q(n2470) );
  AO22X1 U556 ( .IN1(\ram[200][3] ), .IN2(n167), .IN3(n714), .IN4(datain[3]), 
        .Q(n2471) );
  AO22X1 U557 ( .IN1(\ram[200][4] ), .IN2(n167), .IN3(n714), .IN4(datain[4]), 
        .Q(n2472) );
  AO22X1 U558 ( .IN1(\ram[200][5] ), .IN2(n167), .IN3(n714), .IN4(datain[5]), 
        .Q(n2473) );
  AO22X1 U559 ( .IN1(\ram[200][6] ), .IN2(n167), .IN3(n714), .IN4(datain[6]), 
        .Q(n2474) );
  AO22X1 U560 ( .IN1(\ram[200][7] ), .IN2(n167), .IN3(n714), .IN4(datain[7]), 
        .Q(n2475) );
  AO22X1 U563 ( .IN1(\ram[199][0] ), .IN2(n170), .IN3(n567), .IN4(datain[0]), 
        .Q(n2476) );
  AO22X1 U564 ( .IN1(\ram[199][1] ), .IN2(n170), .IN3(n567), .IN4(datain[1]), 
        .Q(n2477) );
  AO22X1 U565 ( .IN1(\ram[199][2] ), .IN2(n170), .IN3(n567), .IN4(datain[2]), 
        .Q(n2478) );
  AO22X1 U566 ( .IN1(\ram[199][3] ), .IN2(n170), .IN3(n567), .IN4(datain[3]), 
        .Q(n2479) );
  AO22X1 U567 ( .IN1(\ram[199][4] ), .IN2(n170), .IN3(n567), .IN4(datain[4]), 
        .Q(n2480) );
  AO22X1 U568 ( .IN1(\ram[199][5] ), .IN2(n170), .IN3(n567), .IN4(datain[5]), 
        .Q(n2481) );
  AO22X1 U569 ( .IN1(\ram[199][6] ), .IN2(n170), .IN3(n567), .IN4(datain[6]), 
        .Q(n2482) );
  AO22X1 U570 ( .IN1(\ram[199][7] ), .IN2(n170), .IN3(n567), .IN4(datain[7]), 
        .Q(n2483) );
  AO22X1 U573 ( .IN1(\ram[198][0] ), .IN2(n173), .IN3(n4160), .IN4(datain[0]), 
        .Q(n2484) );
  AO22X1 U574 ( .IN1(\ram[198][1] ), .IN2(n173), .IN3(n4160), .IN4(datain[1]), 
        .Q(n2485) );
  AO22X1 U575 ( .IN1(\ram[198][2] ), .IN2(n173), .IN3(n4160), .IN4(datain[2]), 
        .Q(n2486) );
  AO22X1 U576 ( .IN1(\ram[198][3] ), .IN2(n173), .IN3(n4160), .IN4(datain[3]), 
        .Q(n2487) );
  AO22X1 U577 ( .IN1(\ram[198][4] ), .IN2(n173), .IN3(n4160), .IN4(datain[4]), 
        .Q(n2488) );
  AO22X1 U578 ( .IN1(\ram[198][5] ), .IN2(n173), .IN3(n4160), .IN4(datain[5]), 
        .Q(n2489) );
  AO22X1 U579 ( .IN1(\ram[198][6] ), .IN2(n173), .IN3(n4160), .IN4(datain[6]), 
        .Q(n2490) );
  AO22X1 U580 ( .IN1(\ram[198][7] ), .IN2(n173), .IN3(n4160), .IN4(datain[7]), 
        .Q(n2491) );
  AO22X1 U583 ( .IN1(\ram[197][0] ), .IN2(n176), .IN3(n663), .IN4(datain[0]), 
        .Q(n2492) );
  AO22X1 U584 ( .IN1(\ram[197][1] ), .IN2(n176), .IN3(n663), .IN4(datain[1]), 
        .Q(n2493) );
  AO22X1 U585 ( .IN1(\ram[197][2] ), .IN2(n176), .IN3(n663), .IN4(datain[2]), 
        .Q(n2494) );
  AO22X1 U586 ( .IN1(\ram[197][3] ), .IN2(n176), .IN3(n663), .IN4(datain[3]), 
        .Q(n2495) );
  AO22X1 U587 ( .IN1(\ram[197][4] ), .IN2(n176), .IN3(n663), .IN4(datain[4]), 
        .Q(n2496) );
  AO22X1 U588 ( .IN1(\ram[197][5] ), .IN2(n176), .IN3(n663), .IN4(datain[5]), 
        .Q(n2497) );
  AO22X1 U589 ( .IN1(\ram[197][6] ), .IN2(n176), .IN3(n663), .IN4(datain[6]), 
        .Q(n2498) );
  AO22X1 U590 ( .IN1(\ram[197][7] ), .IN2(n176), .IN3(n663), .IN4(datain[7]), 
        .Q(n2499) );
  AO22X1 U593 ( .IN1(\ram[196][0] ), .IN2(n179), .IN3(n4112), .IN4(datain[0]), 
        .Q(n2500) );
  AO22X1 U594 ( .IN1(\ram[196][1] ), .IN2(n179), .IN3(n4112), .IN4(datain[1]), 
        .Q(n2501) );
  AO22X1 U595 ( .IN1(\ram[196][2] ), .IN2(n179), .IN3(n4112), .IN4(datain[2]), 
        .Q(n2502) );
  AO22X1 U596 ( .IN1(\ram[196][3] ), .IN2(n179), .IN3(n4112), .IN4(datain[3]), 
        .Q(n2503) );
  AO22X1 U597 ( .IN1(\ram[196][4] ), .IN2(n179), .IN3(n4112), .IN4(datain[4]), 
        .Q(n2504) );
  AO22X1 U598 ( .IN1(\ram[196][5] ), .IN2(n179), .IN3(n4112), .IN4(datain[5]), 
        .Q(n2505) );
  AO22X1 U599 ( .IN1(\ram[196][6] ), .IN2(n179), .IN3(n4112), .IN4(datain[6]), 
        .Q(n2506) );
  AO22X1 U600 ( .IN1(\ram[196][7] ), .IN2(n179), .IN3(n4112), .IN4(datain[7]), 
        .Q(n2507) );
  AO22X1 U603 ( .IN1(\ram[195][0] ), .IN2(n182), .IN3(n519), .IN4(datain[0]), 
        .Q(n2508) );
  AO22X1 U604 ( .IN1(\ram[195][1] ), .IN2(n182), .IN3(n519), .IN4(datain[1]), 
        .Q(n2509) );
  AO22X1 U605 ( .IN1(\ram[195][2] ), .IN2(n182), .IN3(n519), .IN4(datain[2]), 
        .Q(n2510) );
  AO22X1 U606 ( .IN1(\ram[195][3] ), .IN2(n182), .IN3(n519), .IN4(datain[3]), 
        .Q(n2511) );
  AO22X1 U607 ( .IN1(\ram[195][4] ), .IN2(n182), .IN3(n519), .IN4(datain[4]), 
        .Q(n2512) );
  AO22X1 U608 ( .IN1(\ram[195][5] ), .IN2(n182), .IN3(n519), .IN4(datain[5]), 
        .Q(n2513) );
  AO22X1 U609 ( .IN1(\ram[195][6] ), .IN2(n182), .IN3(n519), .IN4(datain[6]), 
        .Q(n2514) );
  AO22X1 U610 ( .IN1(\ram[195][7] ), .IN2(n182), .IN3(n519), .IN4(datain[7]), 
        .Q(n2515) );
  AO22X1 U613 ( .IN1(\ram[194][0] ), .IN2(n185), .IN3(n4143), .IN4(datain[0]), 
        .Q(n2516) );
  AO22X1 U614 ( .IN1(\ram[194][1] ), .IN2(n185), .IN3(n4143), .IN4(datain[1]), 
        .Q(n2517) );
  AO22X1 U615 ( .IN1(\ram[194][2] ), .IN2(n185), .IN3(n4143), .IN4(datain[2]), 
        .Q(n2518) );
  AO22X1 U616 ( .IN1(\ram[194][3] ), .IN2(n185), .IN3(n4143), .IN4(datain[3]), 
        .Q(n2519) );
  AO22X1 U617 ( .IN1(\ram[194][4] ), .IN2(n185), .IN3(n4143), .IN4(datain[4]), 
        .Q(n2520) );
  AO22X1 U618 ( .IN1(\ram[194][5] ), .IN2(n185), .IN3(n4143), .IN4(datain[5]), 
        .Q(n2521) );
  AO22X1 U619 ( .IN1(\ram[194][6] ), .IN2(n185), .IN3(n4143), .IN4(datain[6]), 
        .Q(n2522) );
  AO22X1 U620 ( .IN1(\ram[194][7] ), .IN2(n185), .IN3(n4143), .IN4(datain[7]), 
        .Q(n2523) );
  AO22X1 U623 ( .IN1(\ram[193][0] ), .IN2(n188), .IN3(n615), .IN4(datain[0]), 
        .Q(n2524) );
  AO22X1 U624 ( .IN1(\ram[193][1] ), .IN2(n188), .IN3(n615), .IN4(datain[1]), 
        .Q(n2525) );
  AO22X1 U625 ( .IN1(\ram[193][2] ), .IN2(n188), .IN3(n615), .IN4(datain[2]), 
        .Q(n2526) );
  AO22X1 U626 ( .IN1(\ram[193][3] ), .IN2(n188), .IN3(n615), .IN4(datain[3]), 
        .Q(n2527) );
  AO22X1 U627 ( .IN1(\ram[193][4] ), .IN2(n188), .IN3(n615), .IN4(datain[4]), 
        .Q(n2528) );
  AO22X1 U628 ( .IN1(\ram[193][5] ), .IN2(n188), .IN3(n615), .IN4(datain[5]), 
        .Q(n2529) );
  AO22X1 U629 ( .IN1(\ram[193][6] ), .IN2(n188), .IN3(n615), .IN4(datain[6]), 
        .Q(n2530) );
  AO22X1 U630 ( .IN1(\ram[193][7] ), .IN2(n188), .IN3(n615), .IN4(datain[7]), 
        .Q(n2531) );
  AO22X1 U633 ( .IN1(\ram[192][0] ), .IN2(n191), .IN3(n4134), .IN4(datain[0]), 
        .Q(n2532) );
  AO22X1 U634 ( .IN1(\ram[192][1] ), .IN2(n191), .IN3(n4134), .IN4(datain[1]), 
        .Q(n2533) );
  AO22X1 U635 ( .IN1(\ram[192][2] ), .IN2(n191), .IN3(n4134), .IN4(datain[2]), 
        .Q(n2534) );
  AO22X1 U636 ( .IN1(\ram[192][3] ), .IN2(n191), .IN3(n4134), .IN4(datain[3]), 
        .Q(n2535) );
  AO22X1 U637 ( .IN1(\ram[192][4] ), .IN2(n191), .IN3(n4134), .IN4(datain[4]), 
        .Q(n2536) );
  AO22X1 U638 ( .IN1(\ram[192][5] ), .IN2(n191), .IN3(n4134), .IN4(datain[5]), 
        .Q(n2537) );
  AO22X1 U639 ( .IN1(\ram[192][6] ), .IN2(n191), .IN3(n4134), .IN4(datain[6]), 
        .Q(n2538) );
  AO22X1 U640 ( .IN1(\ram[192][7] ), .IN2(n191), .IN3(n4134), .IN4(datain[7]), 
        .Q(n2539) );
  AO22X1 U643 ( .IN1(\ram[191][0] ), .IN2(n194), .IN3(n393), .IN4(datain[0]), 
        .Q(n2540) );
  AO22X1 U644 ( .IN1(\ram[191][1] ), .IN2(n194), .IN3(n393), .IN4(datain[1]), 
        .Q(n2541) );
  AO22X1 U645 ( .IN1(\ram[191][2] ), .IN2(n194), .IN3(n393), .IN4(datain[2]), 
        .Q(n2542) );
  AO22X1 U646 ( .IN1(\ram[191][3] ), .IN2(n194), .IN3(n393), .IN4(datain[3]), 
        .Q(n2543) );
  AO22X1 U647 ( .IN1(\ram[191][4] ), .IN2(n194), .IN3(n393), .IN4(datain[4]), 
        .Q(n2544) );
  AO22X1 U648 ( .IN1(\ram[191][5] ), .IN2(n194), .IN3(n393), .IN4(datain[5]), 
        .Q(n2545) );
  AO22X1 U649 ( .IN1(\ram[191][6] ), .IN2(n194), .IN3(n393), .IN4(datain[6]), 
        .Q(n2546) );
  AO22X1 U650 ( .IN1(\ram[191][7] ), .IN2(n194), .IN3(n393), .IN4(datain[7]), 
        .Q(n2547) );
  AO22X1 U653 ( .IN1(\ram[190][0] ), .IN2(n197), .IN3(n4089), .IN4(datain[0]), 
        .Q(n2548) );
  AO22X1 U654 ( .IN1(\ram[190][1] ), .IN2(n197), .IN3(n4089), .IN4(datain[1]), 
        .Q(n2549) );
  AO22X1 U655 ( .IN1(\ram[190][2] ), .IN2(n197), .IN3(n4089), .IN4(datain[2]), 
        .Q(n2550) );
  AO22X1 U656 ( .IN1(\ram[190][3] ), .IN2(n197), .IN3(n4089), .IN4(datain[3]), 
        .Q(n2551) );
  AO22X1 U657 ( .IN1(\ram[190][4] ), .IN2(n197), .IN3(n4089), .IN4(datain[4]), 
        .Q(n2552) );
  AO22X1 U658 ( .IN1(\ram[190][5] ), .IN2(n197), .IN3(n4089), .IN4(datain[5]), 
        .Q(n2553) );
  AO22X1 U659 ( .IN1(\ram[190][6] ), .IN2(n197), .IN3(n4089), .IN4(datain[6]), 
        .Q(n2554) );
  AO22X1 U660 ( .IN1(\ram[190][7] ), .IN2(n197), .IN3(n4089), .IN4(datain[7]), 
        .Q(n2555) );
  AO22X1 U663 ( .IN1(\ram[189][0] ), .IN2(n200), .IN3(n450), .IN4(datain[0]), 
        .Q(n2556) );
  AO22X1 U664 ( .IN1(\ram[189][1] ), .IN2(n200), .IN3(n450), .IN4(datain[1]), 
        .Q(n2557) );
  AO22X1 U665 ( .IN1(\ram[189][2] ), .IN2(n200), .IN3(n450), .IN4(datain[2]), 
        .Q(n2558) );
  AO22X1 U666 ( .IN1(\ram[189][3] ), .IN2(n200), .IN3(n450), .IN4(datain[3]), 
        .Q(n2559) );
  AO22X1 U667 ( .IN1(\ram[189][4] ), .IN2(n200), .IN3(n450), .IN4(datain[4]), 
        .Q(n2560) );
  AO22X1 U668 ( .IN1(\ram[189][5] ), .IN2(n200), .IN3(n450), .IN4(datain[5]), 
        .Q(n2561) );
  AO22X1 U669 ( .IN1(\ram[189][6] ), .IN2(n200), .IN3(n450), .IN4(datain[6]), 
        .Q(n2562) );
  AO22X1 U670 ( .IN1(\ram[189][7] ), .IN2(n200), .IN3(n450), .IN4(datain[7]), 
        .Q(n2563) );
  AO22X1 U673 ( .IN1(\ram[188][0] ), .IN2(n203), .IN3(n1974), .IN4(datain[0]), 
        .Q(n2564) );
  AO22X1 U674 ( .IN1(\ram[188][1] ), .IN2(n203), .IN3(n1974), .IN4(datain[1]), 
        .Q(n2565) );
  AO22X1 U675 ( .IN1(\ram[188][2] ), .IN2(n203), .IN3(n1974), .IN4(datain[2]), 
        .Q(n2566) );
  AO22X1 U676 ( .IN1(\ram[188][3] ), .IN2(n203), .IN3(n1974), .IN4(datain[3]), 
        .Q(n2567) );
  AO22X1 U677 ( .IN1(\ram[188][4] ), .IN2(n203), .IN3(n1974), .IN4(datain[4]), 
        .Q(n2568) );
  AO22X1 U678 ( .IN1(\ram[188][5] ), .IN2(n203), .IN3(n1974), .IN4(datain[5]), 
        .Q(n2569) );
  AO22X1 U679 ( .IN1(\ram[188][6] ), .IN2(n203), .IN3(n1974), .IN4(datain[6]), 
        .Q(n2570) );
  AO22X1 U680 ( .IN1(\ram[188][7] ), .IN2(n203), .IN3(n1974), .IN4(datain[7]), 
        .Q(n2571) );
  AO22X1 U683 ( .IN1(\ram[187][0] ), .IN2(n206), .IN3(n339), .IN4(datain[0]), 
        .Q(n2572) );
  AO22X1 U684 ( .IN1(\ram[187][1] ), .IN2(n206), .IN3(n339), .IN4(datain[1]), 
        .Q(n2573) );
  AO22X1 U685 ( .IN1(\ram[187][2] ), .IN2(n206), .IN3(n339), .IN4(datain[2]), 
        .Q(n2574) );
  AO22X1 U686 ( .IN1(\ram[187][3] ), .IN2(n206), .IN3(n339), .IN4(datain[3]), 
        .Q(n2575) );
  AO22X1 U687 ( .IN1(\ram[187][4] ), .IN2(n206), .IN3(n339), .IN4(datain[4]), 
        .Q(n2576) );
  AO22X1 U688 ( .IN1(\ram[187][5] ), .IN2(n206), .IN3(n339), .IN4(datain[5]), 
        .Q(n2577) );
  AO22X1 U689 ( .IN1(\ram[187][6] ), .IN2(n206), .IN3(n339), .IN4(datain[6]), 
        .Q(n2578) );
  AO22X1 U690 ( .IN1(\ram[187][7] ), .IN2(n206), .IN3(n339), .IN4(datain[7]), 
        .Q(n2579) );
  AO22X1 U693 ( .IN1(\ram[186][0] ), .IN2(n209), .IN3(n4085), .IN4(datain[0]), 
        .Q(n2580) );
  AO22X1 U694 ( .IN1(\ram[186][1] ), .IN2(n209), .IN3(n4085), .IN4(datain[1]), 
        .Q(n2581) );
  AO22X1 U695 ( .IN1(\ram[186][2] ), .IN2(n209), .IN3(n4085), .IN4(datain[2]), 
        .Q(n2582) );
  AO22X1 U696 ( .IN1(\ram[186][3] ), .IN2(n209), .IN3(n4085), .IN4(datain[3]), 
        .Q(n2583) );
  AO22X1 U697 ( .IN1(\ram[186][4] ), .IN2(n209), .IN3(n4085), .IN4(datain[4]), 
        .Q(n2584) );
  AO22X1 U698 ( .IN1(\ram[186][5] ), .IN2(n209), .IN3(n4085), .IN4(datain[5]), 
        .Q(n2585) );
  AO22X1 U699 ( .IN1(\ram[186][6] ), .IN2(n209), .IN3(n4085), .IN4(datain[6]), 
        .Q(n2586) );
  AO22X1 U700 ( .IN1(\ram[186][7] ), .IN2(n209), .IN3(n4085), .IN4(datain[7]), 
        .Q(n2587) );
  AO22X1 U703 ( .IN1(\ram[185][0] ), .IN2(n212), .IN3(n438), .IN4(datain[0]), 
        .Q(n2588) );
  AO22X1 U704 ( .IN1(\ram[185][1] ), .IN2(n212), .IN3(n438), .IN4(datain[1]), 
        .Q(n2589) );
  AO22X1 U705 ( .IN1(\ram[185][2] ), .IN2(n212), .IN3(n438), .IN4(datain[2]), 
        .Q(n2590) );
  AO22X1 U706 ( .IN1(\ram[185][3] ), .IN2(n212), .IN3(n438), .IN4(datain[3]), 
        .Q(n2591) );
  AO22X1 U707 ( .IN1(\ram[185][4] ), .IN2(n212), .IN3(n438), .IN4(datain[4]), 
        .Q(n2592) );
  AO22X1 U708 ( .IN1(\ram[185][5] ), .IN2(n212), .IN3(n438), .IN4(datain[5]), 
        .Q(n2593) );
  AO22X1 U709 ( .IN1(\ram[185][6] ), .IN2(n212), .IN3(n438), .IN4(datain[6]), 
        .Q(n2594) );
  AO22X1 U710 ( .IN1(\ram[185][7] ), .IN2(n212), .IN3(n438), .IN4(datain[7]), 
        .Q(n2595) );
  AO22X1 U713 ( .IN1(\ram[184][0] ), .IN2(n215), .IN3(n729), .IN4(datain[0]), 
        .Q(n2596) );
  AO22X1 U714 ( .IN1(\ram[184][1] ), .IN2(n215), .IN3(n729), .IN4(datain[1]), 
        .Q(n2597) );
  AO22X1 U715 ( .IN1(\ram[184][2] ), .IN2(n215), .IN3(n729), .IN4(datain[2]), 
        .Q(n2598) );
  AO22X1 U716 ( .IN1(\ram[184][3] ), .IN2(n215), .IN3(n729), .IN4(datain[3]), 
        .Q(n2599) );
  AO22X1 U717 ( .IN1(\ram[184][4] ), .IN2(n215), .IN3(n729), .IN4(datain[4]), 
        .Q(n2600) );
  AO22X1 U718 ( .IN1(\ram[184][5] ), .IN2(n215), .IN3(n729), .IN4(datain[5]), 
        .Q(n2601) );
  AO22X1 U719 ( .IN1(\ram[184][6] ), .IN2(n215), .IN3(n729), .IN4(datain[6]), 
        .Q(n2602) );
  AO22X1 U720 ( .IN1(\ram[184][7] ), .IN2(n215), .IN3(n729), .IN4(datain[7]), 
        .Q(n2603) );
  AO22X1 U723 ( .IN1(\ram[183][0] ), .IN2(n218), .IN3(n582), .IN4(datain[0]), 
        .Q(n2604) );
  AO22X1 U724 ( .IN1(\ram[183][1] ), .IN2(n218), .IN3(n582), .IN4(datain[1]), 
        .Q(n2605) );
  AO22X1 U725 ( .IN1(\ram[183][2] ), .IN2(n218), .IN3(n582), .IN4(datain[2]), 
        .Q(n2606) );
  AO22X1 U726 ( .IN1(\ram[183][3] ), .IN2(n218), .IN3(n582), .IN4(datain[3]), 
        .Q(n2607) );
  AO22X1 U727 ( .IN1(\ram[183][4] ), .IN2(n218), .IN3(n582), .IN4(datain[4]), 
        .Q(n2608) );
  AO22X1 U728 ( .IN1(\ram[183][5] ), .IN2(n218), .IN3(n582), .IN4(datain[5]), 
        .Q(n2609) );
  AO22X1 U729 ( .IN1(\ram[183][6] ), .IN2(n218), .IN3(n582), .IN4(datain[6]), 
        .Q(n2610) );
  AO22X1 U730 ( .IN1(\ram[183][7] ), .IN2(n218), .IN3(n582), .IN4(datain[7]), 
        .Q(n2611) );
  AO22X1 U733 ( .IN1(\ram[182][0] ), .IN2(n221), .IN3(n4165), .IN4(datain[0]), 
        .Q(n2612) );
  AO22X1 U734 ( .IN1(\ram[182][1] ), .IN2(n221), .IN3(n4165), .IN4(datain[1]), 
        .Q(n2613) );
  AO22X1 U735 ( .IN1(\ram[182][2] ), .IN2(n221), .IN3(n4165), .IN4(datain[2]), 
        .Q(n2614) );
  AO22X1 U736 ( .IN1(\ram[182][3] ), .IN2(n221), .IN3(n4165), .IN4(datain[3]), 
        .Q(n2615) );
  AO22X1 U737 ( .IN1(\ram[182][4] ), .IN2(n221), .IN3(n4165), .IN4(datain[4]), 
        .Q(n2616) );
  AO22X1 U738 ( .IN1(\ram[182][5] ), .IN2(n221), .IN3(n4165), .IN4(datain[5]), 
        .Q(n2617) );
  AO22X1 U739 ( .IN1(\ram[182][6] ), .IN2(n221), .IN3(n4165), .IN4(datain[6]), 
        .Q(n2618) );
  AO22X1 U740 ( .IN1(\ram[182][7] ), .IN2(n221), .IN3(n4165), .IN4(datain[7]), 
        .Q(n2619) );
  AO22X1 U743 ( .IN1(\ram[181][0] ), .IN2(n224), .IN3(n678), .IN4(datain[0]), 
        .Q(n2620) );
  AO22X1 U744 ( .IN1(\ram[181][1] ), .IN2(n224), .IN3(n678), .IN4(datain[1]), 
        .Q(n2621) );
  AO22X1 U745 ( .IN1(\ram[181][2] ), .IN2(n224), .IN3(n678), .IN4(datain[2]), 
        .Q(n2622) );
  AO22X1 U746 ( .IN1(\ram[181][3] ), .IN2(n224), .IN3(n678), .IN4(datain[3]), 
        .Q(n2623) );
  AO22X1 U747 ( .IN1(\ram[181][4] ), .IN2(n224), .IN3(n678), .IN4(datain[4]), 
        .Q(n2624) );
  AO22X1 U748 ( .IN1(\ram[181][5] ), .IN2(n224), .IN3(n678), .IN4(datain[5]), 
        .Q(n2625) );
  AO22X1 U749 ( .IN1(\ram[181][6] ), .IN2(n224), .IN3(n678), .IN4(datain[6]), 
        .Q(n2626) );
  AO22X1 U750 ( .IN1(\ram[181][7] ), .IN2(n224), .IN3(n678), .IN4(datain[7]), 
        .Q(n2627) );
  AO22X1 U753 ( .IN1(\ram[180][0] ), .IN2(n227), .IN3(n4117), .IN4(datain[0]), 
        .Q(n2628) );
  AO22X1 U754 ( .IN1(\ram[180][1] ), .IN2(n227), .IN3(n4117), .IN4(datain[1]), 
        .Q(n2629) );
  AO22X1 U755 ( .IN1(\ram[180][2] ), .IN2(n227), .IN3(n4117), .IN4(datain[2]), 
        .Q(n2630) );
  AO22X1 U756 ( .IN1(\ram[180][3] ), .IN2(n227), .IN3(n4117), .IN4(datain[3]), 
        .Q(n2631) );
  AO22X1 U757 ( .IN1(\ram[180][4] ), .IN2(n227), .IN3(n4117), .IN4(datain[4]), 
        .Q(n2632) );
  AO22X1 U758 ( .IN1(\ram[180][5] ), .IN2(n227), .IN3(n4117), .IN4(datain[5]), 
        .Q(n2633) );
  AO22X1 U759 ( .IN1(\ram[180][6] ), .IN2(n227), .IN3(n4117), .IN4(datain[6]), 
        .Q(n2634) );
  AO22X1 U760 ( .IN1(\ram[180][7] ), .IN2(n227), .IN3(n4117), .IN4(datain[7]), 
        .Q(n2635) );
  AO22X1 U763 ( .IN1(\ram[179][0] ), .IN2(n230), .IN3(n534), .IN4(datain[0]), 
        .Q(n2636) );
  AO22X1 U764 ( .IN1(\ram[179][1] ), .IN2(n230), .IN3(n534), .IN4(datain[1]), 
        .Q(n2637) );
  AO22X1 U765 ( .IN1(\ram[179][2] ), .IN2(n230), .IN3(n534), .IN4(datain[2]), 
        .Q(n2638) );
  AO22X1 U766 ( .IN1(\ram[179][3] ), .IN2(n230), .IN3(n534), .IN4(datain[3]), 
        .Q(n2639) );
  AO22X1 U767 ( .IN1(\ram[179][4] ), .IN2(n230), .IN3(n534), .IN4(datain[4]), 
        .Q(n2640) );
  AO22X1 U768 ( .IN1(\ram[179][5] ), .IN2(n230), .IN3(n534), .IN4(datain[5]), 
        .Q(n2641) );
  AO22X1 U769 ( .IN1(\ram[179][6] ), .IN2(n230), .IN3(n534), .IN4(datain[6]), 
        .Q(n2642) );
  AO22X1 U770 ( .IN1(\ram[179][7] ), .IN2(n230), .IN3(n534), .IN4(datain[7]), 
        .Q(n2643) );
  AO22X1 U773 ( .IN1(\ram[178][0] ), .IN2(n233), .IN3(n4149), .IN4(datain[0]), 
        .Q(n2644) );
  AO22X1 U774 ( .IN1(\ram[178][1] ), .IN2(n233), .IN3(n4149), .IN4(datain[1]), 
        .Q(n2645) );
  AO22X1 U775 ( .IN1(\ram[178][2] ), .IN2(n233), .IN3(n4149), .IN4(datain[2]), 
        .Q(n2646) );
  AO22X1 U776 ( .IN1(\ram[178][3] ), .IN2(n233), .IN3(n4149), .IN4(datain[3]), 
        .Q(n2647) );
  AO22X1 U777 ( .IN1(\ram[178][4] ), .IN2(n233), .IN3(n4149), .IN4(datain[4]), 
        .Q(n2648) );
  AO22X1 U778 ( .IN1(\ram[178][5] ), .IN2(n233), .IN3(n4149), .IN4(datain[5]), 
        .Q(n2649) );
  AO22X1 U779 ( .IN1(\ram[178][6] ), .IN2(n233), .IN3(n4149), .IN4(datain[6]), 
        .Q(n2650) );
  AO22X1 U780 ( .IN1(\ram[178][7] ), .IN2(n233), .IN3(n4149), .IN4(datain[7]), 
        .Q(n2651) );
  AO22X1 U783 ( .IN1(\ram[177][0] ), .IN2(n236), .IN3(n630), .IN4(datain[0]), 
        .Q(n2652) );
  AO22X1 U784 ( .IN1(\ram[177][1] ), .IN2(n236), .IN3(n630), .IN4(datain[1]), 
        .Q(n2653) );
  AO22X1 U785 ( .IN1(\ram[177][2] ), .IN2(n236), .IN3(n630), .IN4(datain[2]), 
        .Q(n2654) );
  AO22X1 U786 ( .IN1(\ram[177][3] ), .IN2(n236), .IN3(n630), .IN4(datain[3]), 
        .Q(n2655) );
  AO22X1 U787 ( .IN1(\ram[177][4] ), .IN2(n236), .IN3(n630), .IN4(datain[4]), 
        .Q(n2656) );
  AO22X1 U788 ( .IN1(\ram[177][5] ), .IN2(n236), .IN3(n630), .IN4(datain[5]), 
        .Q(n2657) );
  AO22X1 U789 ( .IN1(\ram[177][6] ), .IN2(n236), .IN3(n630), .IN4(datain[6]), 
        .Q(n2658) );
  AO22X1 U790 ( .IN1(\ram[177][7] ), .IN2(n236), .IN3(n630), .IN4(datain[7]), 
        .Q(n2659) );
  AO22X1 U793 ( .IN1(\ram[176][0] ), .IN2(n239), .IN3(n4131), .IN4(datain[0]), 
        .Q(n2660) );
  AO22X1 U794 ( .IN1(\ram[176][1] ), .IN2(n239), .IN3(n4131), .IN4(datain[1]), 
        .Q(n2661) );
  AO22X1 U795 ( .IN1(\ram[176][2] ), .IN2(n239), .IN3(n4131), .IN4(datain[2]), 
        .Q(n2662) );
  AO22X1 U796 ( .IN1(\ram[176][3] ), .IN2(n239), .IN3(n4131), .IN4(datain[3]), 
        .Q(n2663) );
  AO22X1 U797 ( .IN1(\ram[176][4] ), .IN2(n239), .IN3(n4131), .IN4(datain[4]), 
        .Q(n2664) );
  AO22X1 U798 ( .IN1(\ram[176][5] ), .IN2(n239), .IN3(n4131), .IN4(datain[5]), 
        .Q(n2665) );
  AO22X1 U799 ( .IN1(\ram[176][6] ), .IN2(n239), .IN3(n4131), .IN4(datain[6]), 
        .Q(n2666) );
  AO22X1 U800 ( .IN1(\ram[176][7] ), .IN2(n239), .IN3(n4131), .IN4(datain[7]), 
        .Q(n2667) );
  AO22X1 U803 ( .IN1(\ram[175][0] ), .IN2(n242), .IN3(n384), .IN4(datain[0]), 
        .Q(n2668) );
  AO22X1 U804 ( .IN1(\ram[175][1] ), .IN2(n242), .IN3(n384), .IN4(datain[1]), 
        .Q(n2669) );
  AO22X1 U805 ( .IN1(\ram[175][2] ), .IN2(n242), .IN3(n384), .IN4(datain[2]), 
        .Q(n2670) );
  AO22X1 U806 ( .IN1(\ram[175][3] ), .IN2(n242), .IN3(n384), .IN4(datain[3]), 
        .Q(n2671) );
  AO22X1 U807 ( .IN1(\ram[175][4] ), .IN2(n242), .IN3(n384), .IN4(datain[4]), 
        .Q(n2672) );
  AO22X1 U808 ( .IN1(\ram[175][5] ), .IN2(n242), .IN3(n384), .IN4(datain[5]), 
        .Q(n2673) );
  AO22X1 U809 ( .IN1(\ram[175][6] ), .IN2(n242), .IN3(n384), .IN4(datain[6]), 
        .Q(n2674) );
  AO22X1 U810 ( .IN1(\ram[175][7] ), .IN2(n242), .IN3(n384), .IN4(datain[7]), 
        .Q(n2675) );
  AO22X1 U813 ( .IN1(\ram[174][0] ), .IN2(n245), .IN3(n4102), .IN4(datain[0]), 
        .Q(n2676) );
  AO22X1 U814 ( .IN1(\ram[174][1] ), .IN2(n245), .IN3(n4102), .IN4(datain[1]), 
        .Q(n2677) );
  AO22X1 U815 ( .IN1(\ram[174][2] ), .IN2(n245), .IN3(n4102), .IN4(datain[2]), 
        .Q(n2678) );
  AO22X1 U816 ( .IN1(\ram[174][3] ), .IN2(n245), .IN3(n4102), .IN4(datain[3]), 
        .Q(n2679) );
  AO22X1 U817 ( .IN1(\ram[174][4] ), .IN2(n245), .IN3(n4102), .IN4(datain[4]), 
        .Q(n2680) );
  AO22X1 U818 ( .IN1(\ram[174][5] ), .IN2(n245), .IN3(n4102), .IN4(datain[5]), 
        .Q(n2681) );
  AO22X1 U819 ( .IN1(\ram[174][6] ), .IN2(n245), .IN3(n4102), .IN4(datain[6]), 
        .Q(n2682) );
  AO22X1 U820 ( .IN1(\ram[174][7] ), .IN2(n245), .IN3(n4102), .IN4(datain[7]), 
        .Q(n2683) );
  AO22X1 U823 ( .IN1(\ram[173][0] ), .IN2(n248), .IN3(n489), .IN4(datain[0]), 
        .Q(n2684) );
  AO22X1 U824 ( .IN1(\ram[173][1] ), .IN2(n248), .IN3(n489), .IN4(datain[1]), 
        .Q(n2685) );
  AO22X1 U825 ( .IN1(\ram[173][2] ), .IN2(n248), .IN3(n489), .IN4(datain[2]), 
        .Q(n2686) );
  AO22X1 U826 ( .IN1(\ram[173][3] ), .IN2(n248), .IN3(n489), .IN4(datain[3]), 
        .Q(n2687) );
  AO22X1 U827 ( .IN1(\ram[173][4] ), .IN2(n248), .IN3(n489), .IN4(datain[4]), 
        .Q(n2688) );
  AO22X1 U828 ( .IN1(\ram[173][5] ), .IN2(n248), .IN3(n489), .IN4(datain[5]), 
        .Q(n2689) );
  AO22X1 U829 ( .IN1(\ram[173][6] ), .IN2(n248), .IN3(n489), .IN4(datain[6]), 
        .Q(n2690) );
  AO22X1 U830 ( .IN1(\ram[173][7] ), .IN2(n248), .IN3(n489), .IN4(datain[7]), 
        .Q(n2691) );
  AO22X1 U833 ( .IN1(\ram[172][0] ), .IN2(n251), .IN3(n1975), .IN4(datain[0]), 
        .Q(n2692) );
  AO22X1 U834 ( .IN1(\ram[172][1] ), .IN2(n251), .IN3(n1975), .IN4(datain[1]), 
        .Q(n2693) );
  AO22X1 U835 ( .IN1(\ram[172][2] ), .IN2(n251), .IN3(n1975), .IN4(datain[2]), 
        .Q(n2694) );
  AO22X1 U836 ( .IN1(\ram[172][3] ), .IN2(n251), .IN3(n1975), .IN4(datain[3]), 
        .Q(n2695) );
  AO22X1 U837 ( .IN1(\ram[172][4] ), .IN2(n251), .IN3(n1975), .IN4(datain[4]), 
        .Q(n2696) );
  AO22X1 U838 ( .IN1(\ram[172][5] ), .IN2(n251), .IN3(n1975), .IN4(datain[5]), 
        .Q(n2697) );
  AO22X1 U839 ( .IN1(\ram[172][6] ), .IN2(n251), .IN3(n1975), .IN4(datain[6]), 
        .Q(n2698) );
  AO22X1 U840 ( .IN1(\ram[172][7] ), .IN2(n251), .IN3(n1975), .IN4(datain[7]), 
        .Q(n2699) );
  AO22X1 U843 ( .IN1(\ram[171][0] ), .IN2(n254), .IN3(n342), .IN4(datain[0]), 
        .Q(n2700) );
  AO22X1 U844 ( .IN1(\ram[171][1] ), .IN2(n254), .IN3(n342), .IN4(datain[1]), 
        .Q(n2701) );
  AO22X1 U845 ( .IN1(\ram[171][2] ), .IN2(n254), .IN3(n342), .IN4(datain[2]), 
        .Q(n2702) );
  AO22X1 U846 ( .IN1(\ram[171][3] ), .IN2(n254), .IN3(n342), .IN4(datain[3]), 
        .Q(n2703) );
  AO22X1 U847 ( .IN1(\ram[171][4] ), .IN2(n254), .IN3(n342), .IN4(datain[4]), 
        .Q(n2704) );
  AO22X1 U848 ( .IN1(\ram[171][5] ), .IN2(n254), .IN3(n342), .IN4(datain[5]), 
        .Q(n2705) );
  AO22X1 U849 ( .IN1(\ram[171][6] ), .IN2(n254), .IN3(n342), .IN4(datain[6]), 
        .Q(n2706) );
  AO22X1 U850 ( .IN1(\ram[171][7] ), .IN2(n254), .IN3(n342), .IN4(datain[7]), 
        .Q(n2707) );
  AO22X1 U853 ( .IN1(\ram[170][0] ), .IN2(n257), .IN3(n4086), .IN4(datain[0]), 
        .Q(n2708) );
  AO22X1 U854 ( .IN1(\ram[170][1] ), .IN2(n257), .IN3(n4086), .IN4(datain[1]), 
        .Q(n2709) );
  AO22X1 U855 ( .IN1(\ram[170][2] ), .IN2(n257), .IN3(n4086), .IN4(datain[2]), 
        .Q(n2710) );
  AO22X1 U856 ( .IN1(\ram[170][3] ), .IN2(n257), .IN3(n4086), .IN4(datain[3]), 
        .Q(n2711) );
  AO22X1 U857 ( .IN1(\ram[170][4] ), .IN2(n257), .IN3(n4086), .IN4(datain[4]), 
        .Q(n2712) );
  AO22X1 U858 ( .IN1(\ram[170][5] ), .IN2(n257), .IN3(n4086), .IN4(datain[5]), 
        .Q(n2713) );
  AO22X1 U859 ( .IN1(\ram[170][6] ), .IN2(n257), .IN3(n4086), .IN4(datain[6]), 
        .Q(n2714) );
  AO22X1 U860 ( .IN1(\ram[170][7] ), .IN2(n257), .IN3(n4086), .IN4(datain[7]), 
        .Q(n2715) );
  AO22X1 U863 ( .IN1(\ram[169][0] ), .IN2(n260), .IN3(n441), .IN4(datain[0]), 
        .Q(n2716) );
  AO22X1 U864 ( .IN1(\ram[169][1] ), .IN2(n260), .IN3(n441), .IN4(datain[1]), 
        .Q(n2717) );
  AO22X1 U865 ( .IN1(\ram[169][2] ), .IN2(n260), .IN3(n441), .IN4(datain[2]), 
        .Q(n2718) );
  AO22X1 U866 ( .IN1(\ram[169][3] ), .IN2(n260), .IN3(n441), .IN4(datain[3]), 
        .Q(n2719) );
  AO22X1 U867 ( .IN1(\ram[169][4] ), .IN2(n260), .IN3(n441), .IN4(datain[4]), 
        .Q(n2720) );
  AO22X1 U868 ( .IN1(\ram[169][5] ), .IN2(n260), .IN3(n441), .IN4(datain[5]), 
        .Q(n2721) );
  AO22X1 U869 ( .IN1(\ram[169][6] ), .IN2(n260), .IN3(n441), .IN4(datain[6]), 
        .Q(n2722) );
  AO22X1 U870 ( .IN1(\ram[169][7] ), .IN2(n260), .IN3(n441), .IN4(datain[7]), 
        .Q(n2723) );
  AO22X1 U873 ( .IN1(\ram[168][0] ), .IN2(n263), .IN3(n732), .IN4(datain[0]), 
        .Q(n2724) );
  AO22X1 U874 ( .IN1(\ram[168][1] ), .IN2(n263), .IN3(n732), .IN4(datain[1]), 
        .Q(n2725) );
  AO22X1 U875 ( .IN1(\ram[168][2] ), .IN2(n263), .IN3(n732), .IN4(datain[2]), 
        .Q(n2726) );
  AO22X1 U876 ( .IN1(\ram[168][3] ), .IN2(n263), .IN3(n732), .IN4(datain[3]), 
        .Q(n2727) );
  AO22X1 U877 ( .IN1(\ram[168][4] ), .IN2(n263), .IN3(n732), .IN4(datain[4]), 
        .Q(n2728) );
  AO22X1 U878 ( .IN1(\ram[168][5] ), .IN2(n263), .IN3(n732), .IN4(datain[5]), 
        .Q(n2729) );
  AO22X1 U879 ( .IN1(\ram[168][6] ), .IN2(n263), .IN3(n732), .IN4(datain[6]), 
        .Q(n2730) );
  AO22X1 U880 ( .IN1(\ram[168][7] ), .IN2(n263), .IN3(n732), .IN4(datain[7]), 
        .Q(n2731) );
  AO22X1 U883 ( .IN1(\ram[167][0] ), .IN2(n266), .IN3(n585), .IN4(datain[0]), 
        .Q(n2732) );
  AO22X1 U884 ( .IN1(\ram[167][1] ), .IN2(n266), .IN3(n585), .IN4(datain[1]), 
        .Q(n2733) );
  AO22X1 U885 ( .IN1(\ram[167][2] ), .IN2(n266), .IN3(n585), .IN4(datain[2]), 
        .Q(n2734) );
  AO22X1 U886 ( .IN1(\ram[167][3] ), .IN2(n266), .IN3(n585), .IN4(datain[3]), 
        .Q(n2735) );
  AO22X1 U887 ( .IN1(\ram[167][4] ), .IN2(n266), .IN3(n585), .IN4(datain[4]), 
        .Q(n2736) );
  AO22X1 U888 ( .IN1(\ram[167][5] ), .IN2(n266), .IN3(n585), .IN4(datain[5]), 
        .Q(n2737) );
  AO22X1 U889 ( .IN1(\ram[167][6] ), .IN2(n266), .IN3(n585), .IN4(datain[6]), 
        .Q(n2738) );
  AO22X1 U890 ( .IN1(\ram[167][7] ), .IN2(n266), .IN3(n585), .IN4(datain[7]), 
        .Q(n2739) );
  AO22X1 U893 ( .IN1(\ram[166][0] ), .IN2(n269), .IN3(n4166), .IN4(datain[0]), 
        .Q(n2740) );
  AO22X1 U894 ( .IN1(\ram[166][1] ), .IN2(n269), .IN3(n4166), .IN4(datain[1]), 
        .Q(n2741) );
  AO22X1 U895 ( .IN1(\ram[166][2] ), .IN2(n269), .IN3(n4166), .IN4(datain[2]), 
        .Q(n2742) );
  AO22X1 U896 ( .IN1(\ram[166][3] ), .IN2(n269), .IN3(n4166), .IN4(datain[3]), 
        .Q(n2743) );
  AO22X1 U897 ( .IN1(\ram[166][4] ), .IN2(n269), .IN3(n4166), .IN4(datain[4]), 
        .Q(n2744) );
  AO22X1 U898 ( .IN1(\ram[166][5] ), .IN2(n269), .IN3(n4166), .IN4(datain[5]), 
        .Q(n2745) );
  AO22X1 U899 ( .IN1(\ram[166][6] ), .IN2(n269), .IN3(n4166), .IN4(datain[6]), 
        .Q(n2746) );
  AO22X1 U900 ( .IN1(\ram[166][7] ), .IN2(n269), .IN3(n4166), .IN4(datain[7]), 
        .Q(n2747) );
  AO22X1 U903 ( .IN1(\ram[165][0] ), .IN2(n272), .IN3(n681), .IN4(n63), .Q(
        n2748) );
  AO22X1 U904 ( .IN1(\ram[165][1] ), .IN2(n272), .IN3(n681), .IN4(n96), .Q(
        n2749) );
  AO22X1 U905 ( .IN1(\ram[165][2] ), .IN2(n272), .IN3(n681), .IN4(n129), .Q(
        n2750) );
  AO22X1 U906 ( .IN1(\ram[165][3] ), .IN2(n272), .IN3(n681), .IN4(n162), .Q(
        n2751) );
  AO22X1 U907 ( .IN1(\ram[165][4] ), .IN2(n272), .IN3(n681), .IN4(n195), .Q(
        n2752) );
  AO22X1 U908 ( .IN1(\ram[165][5] ), .IN2(n272), .IN3(n681), .IN4(n228), .Q(
        n2753) );
  AO22X1 U909 ( .IN1(\ram[165][6] ), .IN2(n272), .IN3(n681), .IN4(n261), .Q(
        n2754) );
  AO22X1 U910 ( .IN1(\ram[165][7] ), .IN2(n272), .IN3(n681), .IN4(n294), .Q(
        n2755) );
  AO22X1 U913 ( .IN1(\ram[164][0] ), .IN2(n275), .IN3(n4118), .IN4(datain[0]), 
        .Q(n2756) );
  AO22X1 U914 ( .IN1(\ram[164][1] ), .IN2(n275), .IN3(n4118), .IN4(datain[1]), 
        .Q(n2757) );
  AO22X1 U915 ( .IN1(\ram[164][2] ), .IN2(n275), .IN3(n4118), .IN4(datain[2]), 
        .Q(n2758) );
  AO22X1 U916 ( .IN1(\ram[164][3] ), .IN2(n275), .IN3(n4118), .IN4(datain[3]), 
        .Q(n2759) );
  AO22X1 U917 ( .IN1(\ram[164][4] ), .IN2(n275), .IN3(n4118), .IN4(datain[4]), 
        .Q(n2760) );
  AO22X1 U918 ( .IN1(\ram[164][5] ), .IN2(n275), .IN3(n4118), .IN4(datain[5]), 
        .Q(n2761) );
  AO22X1 U919 ( .IN1(\ram[164][6] ), .IN2(n275), .IN3(n4118), .IN4(datain[6]), 
        .Q(n2762) );
  AO22X1 U920 ( .IN1(\ram[164][7] ), .IN2(n275), .IN3(n4118), .IN4(datain[7]), 
        .Q(n2763) );
  AO22X1 U923 ( .IN1(\ram[163][0] ), .IN2(n278), .IN3(n537), .IN4(datain[0]), 
        .Q(n2764) );
  AO22X1 U924 ( .IN1(\ram[163][1] ), .IN2(n278), .IN3(n537), .IN4(datain[1]), 
        .Q(n2765) );
  AO22X1 U925 ( .IN1(\ram[163][2] ), .IN2(n278), .IN3(n537), .IN4(datain[2]), 
        .Q(n2766) );
  AO22X1 U926 ( .IN1(\ram[163][3] ), .IN2(n278), .IN3(n537), .IN4(datain[3]), 
        .Q(n2767) );
  AO22X1 U927 ( .IN1(\ram[163][4] ), .IN2(n278), .IN3(n537), .IN4(datain[4]), 
        .Q(n2768) );
  AO22X1 U928 ( .IN1(\ram[163][5] ), .IN2(n278), .IN3(n537), .IN4(datain[5]), 
        .Q(n2769) );
  AO22X1 U929 ( .IN1(\ram[163][6] ), .IN2(n278), .IN3(n537), .IN4(datain[6]), 
        .Q(n2770) );
  AO22X1 U930 ( .IN1(\ram[163][7] ), .IN2(n278), .IN3(n537), .IN4(datain[7]), 
        .Q(n2771) );
  AO22X1 U933 ( .IN1(\ram[162][0] ), .IN2(n281), .IN3(n4150), .IN4(datain[0]), 
        .Q(n2772) );
  AO22X1 U934 ( .IN1(\ram[162][1] ), .IN2(n281), .IN3(n4150), .IN4(datain[1]), 
        .Q(n2773) );
  AO22X1 U935 ( .IN1(\ram[162][2] ), .IN2(n281), .IN3(n4150), .IN4(datain[2]), 
        .Q(n2774) );
  AO22X1 U936 ( .IN1(\ram[162][3] ), .IN2(n281), .IN3(n4150), .IN4(datain[3]), 
        .Q(n2775) );
  AO22X1 U937 ( .IN1(\ram[162][4] ), .IN2(n281), .IN3(n4150), .IN4(datain[4]), 
        .Q(n2776) );
  AO22X1 U938 ( .IN1(\ram[162][5] ), .IN2(n281), .IN3(n4150), .IN4(datain[5]), 
        .Q(n2777) );
  AO22X1 U939 ( .IN1(\ram[162][6] ), .IN2(n281), .IN3(n4150), .IN4(datain[6]), 
        .Q(n2778) );
  AO22X1 U940 ( .IN1(\ram[162][7] ), .IN2(n281), .IN3(n4150), .IN4(datain[7]), 
        .Q(n2779) );
  AO22X1 U943 ( .IN1(\ram[161][0] ), .IN2(n284), .IN3(n633), .IN4(datain[0]), 
        .Q(n2780) );
  AO22X1 U944 ( .IN1(\ram[161][1] ), .IN2(n284), .IN3(n633), .IN4(datain[1]), 
        .Q(n2781) );
  AO22X1 U945 ( .IN1(\ram[161][2] ), .IN2(n284), .IN3(n633), .IN4(datain[2]), 
        .Q(n2782) );
  AO22X1 U946 ( .IN1(\ram[161][3] ), .IN2(n284), .IN3(n633), .IN4(datain[3]), 
        .Q(n2783) );
  AO22X1 U947 ( .IN1(\ram[161][4] ), .IN2(n284), .IN3(n633), .IN4(datain[4]), 
        .Q(n2784) );
  AO22X1 U948 ( .IN1(\ram[161][5] ), .IN2(n284), .IN3(n633), .IN4(datain[5]), 
        .Q(n2785) );
  AO22X1 U949 ( .IN1(\ram[161][6] ), .IN2(n284), .IN3(n633), .IN4(datain[6]), 
        .Q(n2786) );
  AO22X1 U950 ( .IN1(\ram[161][7] ), .IN2(n284), .IN3(n633), .IN4(datain[7]), 
        .Q(n2787) );
  AO22X1 U953 ( .IN1(\ram[160][0] ), .IN2(n287), .IN3(n4129), .IN4(datain[0]), 
        .Q(n2788) );
  AO22X1 U954 ( .IN1(\ram[160][1] ), .IN2(n287), .IN3(n4129), .IN4(datain[1]), 
        .Q(n2789) );
  AO22X1 U955 ( .IN1(\ram[160][2] ), .IN2(n287), .IN3(n4129), .IN4(datain[2]), 
        .Q(n2790) );
  AO22X1 U956 ( .IN1(\ram[160][3] ), .IN2(n287), .IN3(n4129), .IN4(datain[3]), 
        .Q(n2791) );
  AO22X1 U957 ( .IN1(\ram[160][4] ), .IN2(n287), .IN3(n4129), .IN4(datain[4]), 
        .Q(n2792) );
  AO22X1 U958 ( .IN1(\ram[160][5] ), .IN2(n287), .IN3(n4129), .IN4(datain[5]), 
        .Q(n2793) );
  AO22X1 U959 ( .IN1(\ram[160][6] ), .IN2(n287), .IN3(n4129), .IN4(datain[6]), 
        .Q(n2794) );
  AO22X1 U960 ( .IN1(\ram[160][7] ), .IN2(n287), .IN3(n4129), .IN4(datain[7]), 
        .Q(n2795) );
  AO22X1 U963 ( .IN1(\ram[159][0] ), .IN2(n290), .IN3(n378), .IN4(datain[0]), 
        .Q(n2796) );
  AO22X1 U964 ( .IN1(\ram[159][1] ), .IN2(n290), .IN3(n378), .IN4(datain[1]), 
        .Q(n2797) );
  AO22X1 U965 ( .IN1(\ram[159][2] ), .IN2(n290), .IN3(n378), .IN4(datain[2]), 
        .Q(n2798) );
  AO22X1 U966 ( .IN1(\ram[159][3] ), .IN2(n290), .IN3(n378), .IN4(datain[3]), 
        .Q(n2799) );
  AO22X1 U967 ( .IN1(\ram[159][4] ), .IN2(n290), .IN3(n378), .IN4(datain[4]), 
        .Q(n2800) );
  AO22X1 U968 ( .IN1(\ram[159][5] ), .IN2(n290), .IN3(n378), .IN4(datain[5]), 
        .Q(n2801) );
  AO22X1 U969 ( .IN1(\ram[159][6] ), .IN2(n290), .IN3(n378), .IN4(datain[6]), 
        .Q(n2802) );
  AO22X1 U970 ( .IN1(\ram[159][7] ), .IN2(n290), .IN3(n378), .IN4(datain[7]), 
        .Q(n2803) );
  AO22X1 U973 ( .IN1(\ram[158][0] ), .IN2(n293), .IN3(n4100), .IN4(datain[0]), 
        .Q(n2804) );
  AO22X1 U974 ( .IN1(\ram[158][1] ), .IN2(n293), .IN3(n4100), .IN4(datain[1]), 
        .Q(n2805) );
  AO22X1 U975 ( .IN1(\ram[158][2] ), .IN2(n293), .IN3(n4100), .IN4(datain[2]), 
        .Q(n2806) );
  AO22X1 U976 ( .IN1(\ram[158][3] ), .IN2(n293), .IN3(n4100), .IN4(datain[3]), 
        .Q(n2807) );
  AO22X1 U977 ( .IN1(\ram[158][4] ), .IN2(n293), .IN3(n4100), .IN4(datain[4]), 
        .Q(n2808) );
  AO22X1 U978 ( .IN1(\ram[158][5] ), .IN2(n293), .IN3(n4100), .IN4(datain[5]), 
        .Q(n2809) );
  AO22X1 U979 ( .IN1(\ram[158][6] ), .IN2(n293), .IN3(n4100), .IN4(datain[6]), 
        .Q(n2810) );
  AO22X1 U980 ( .IN1(\ram[158][7] ), .IN2(n293), .IN3(n4100), .IN4(datain[7]), 
        .Q(n2811) );
  AO22X1 U983 ( .IN1(\ram[157][0] ), .IN2(n296), .IN3(n483), .IN4(datain[0]), 
        .Q(n2812) );
  AO22X1 U984 ( .IN1(\ram[157][1] ), .IN2(n296), .IN3(n483), .IN4(datain[1]), 
        .Q(n2813) );
  AO22X1 U985 ( .IN1(\ram[157][2] ), .IN2(n296), .IN3(n483), .IN4(datain[2]), 
        .Q(n2814) );
  AO22X1 U986 ( .IN1(\ram[157][3] ), .IN2(n296), .IN3(n483), .IN4(datain[3]), 
        .Q(n2815) );
  AO22X1 U987 ( .IN1(\ram[157][4] ), .IN2(n296), .IN3(n483), .IN4(datain[4]), 
        .Q(n2816) );
  AO22X1 U988 ( .IN1(\ram[157][5] ), .IN2(n296), .IN3(n483), .IN4(datain[5]), 
        .Q(n2817) );
  AO22X1 U989 ( .IN1(\ram[157][6] ), .IN2(n296), .IN3(n483), .IN4(datain[6]), 
        .Q(n2818) );
  AO22X1 U990 ( .IN1(\ram[157][7] ), .IN2(n296), .IN3(n483), .IN4(datain[7]), 
        .Q(n2819) );
  AO22X1 U993 ( .IN1(\ram[156][0] ), .IN2(n299), .IN3(n768), .IN4(datain[0]), 
        .Q(n2820) );
  AO22X1 U994 ( .IN1(\ram[156][1] ), .IN2(n299), .IN3(n768), .IN4(datain[1]), 
        .Q(n2821) );
  AO22X1 U995 ( .IN1(\ram[156][2] ), .IN2(n299), .IN3(n768), .IN4(datain[2]), 
        .Q(n2822) );
  AO22X1 U996 ( .IN1(\ram[156][3] ), .IN2(n299), .IN3(n768), .IN4(datain[3]), 
        .Q(n2823) );
  AO22X1 U997 ( .IN1(\ram[156][4] ), .IN2(n299), .IN3(n768), .IN4(datain[4]), 
        .Q(n2824) );
  AO22X1 U998 ( .IN1(\ram[156][5] ), .IN2(n299), .IN3(n768), .IN4(datain[5]), 
        .Q(n2825) );
  AO22X1 U999 ( .IN1(\ram[156][6] ), .IN2(n299), .IN3(n768), .IN4(datain[6]), 
        .Q(n2826) );
  AO22X1 U1000 ( .IN1(\ram[156][7] ), .IN2(n299), .IN3(n768), .IN4(datain[7]), 
        .Q(n2827) );
  AO22X1 U1003 ( .IN1(\ram[155][0] ), .IN2(n302), .IN3(n333), .IN4(datain[0]), 
        .Q(n2828) );
  AO22X1 U1004 ( .IN1(\ram[155][1] ), .IN2(n302), .IN3(n333), .IN4(datain[1]), 
        .Q(n2829) );
  AO22X1 U1005 ( .IN1(\ram[155][2] ), .IN2(n302), .IN3(n333), .IN4(datain[2]), 
        .Q(n2830) );
  AO22X1 U1006 ( .IN1(\ram[155][3] ), .IN2(n302), .IN3(n333), .IN4(datain[3]), 
        .Q(n2831) );
  AO22X1 U1007 ( .IN1(\ram[155][4] ), .IN2(n302), .IN3(n333), .IN4(datain[4]), 
        .Q(n2832) );
  AO22X1 U1008 ( .IN1(\ram[155][5] ), .IN2(n302), .IN3(n333), .IN4(datain[5]), 
        .Q(n2833) );
  AO22X1 U1009 ( .IN1(\ram[155][6] ), .IN2(n302), .IN3(n333), .IN4(datain[6]), 
        .Q(n2834) );
  AO22X1 U1010 ( .IN1(\ram[155][7] ), .IN2(n302), .IN3(n333), .IN4(datain[7]), 
        .Q(n2835) );
  AO22X1 U1013 ( .IN1(\ram[154][0] ), .IN2(n305), .IN3(n4083), .IN4(datain[0]), 
        .Q(n2836) );
  AO22X1 U1014 ( .IN1(\ram[154][1] ), .IN2(n305), .IN3(n4083), .IN4(datain[1]), 
        .Q(n2837) );
  AO22X1 U1015 ( .IN1(\ram[154][2] ), .IN2(n305), .IN3(n4083), .IN4(datain[2]), 
        .Q(n2838) );
  AO22X1 U1016 ( .IN1(\ram[154][3] ), .IN2(n305), .IN3(n4083), .IN4(datain[3]), 
        .Q(n2839) );
  AO22X1 U1017 ( .IN1(\ram[154][4] ), .IN2(n305), .IN3(n4083), .IN4(datain[4]), 
        .Q(n2840) );
  AO22X1 U1018 ( .IN1(\ram[154][5] ), .IN2(n305), .IN3(n4083), .IN4(datain[5]), 
        .Q(n2841) );
  AO22X1 U1019 ( .IN1(\ram[154][6] ), .IN2(n305), .IN3(n4083), .IN4(datain[6]), 
        .Q(n2842) );
  AO22X1 U1020 ( .IN1(\ram[154][7] ), .IN2(n305), .IN3(n4083), .IN4(datain[7]), 
        .Q(n2843) );
  AO22X1 U1023 ( .IN1(\ram[153][0] ), .IN2(n308), .IN3(n432), .IN4(datain[0]), 
        .Q(n2844) );
  AO22X1 U1024 ( .IN1(\ram[153][1] ), .IN2(n308), .IN3(n432), .IN4(datain[1]), 
        .Q(n2845) );
  AO22X1 U1025 ( .IN1(\ram[153][2] ), .IN2(n308), .IN3(n432), .IN4(datain[2]), 
        .Q(n2846) );
  AO22X1 U1026 ( .IN1(\ram[153][3] ), .IN2(n308), .IN3(n432), .IN4(datain[3]), 
        .Q(n2847) );
  AO22X1 U1027 ( .IN1(\ram[153][4] ), .IN2(n308), .IN3(n432), .IN4(datain[4]), 
        .Q(n2848) );
  AO22X1 U1028 ( .IN1(\ram[153][5] ), .IN2(n308), .IN3(n432), .IN4(datain[5]), 
        .Q(n2849) );
  AO22X1 U1029 ( .IN1(\ram[153][6] ), .IN2(n308), .IN3(n432), .IN4(datain[6]), 
        .Q(n2850) );
  AO22X1 U1030 ( .IN1(\ram[153][7] ), .IN2(n308), .IN3(n432), .IN4(datain[7]), 
        .Q(n2851) );
  AO22X1 U1033 ( .IN1(\ram[152][0] ), .IN2(n311), .IN3(n723), .IN4(datain[0]), 
        .Q(n2852) );
  AO22X1 U1034 ( .IN1(\ram[152][1] ), .IN2(n311), .IN3(n723), .IN4(datain[1]), 
        .Q(n2853) );
  AO22X1 U1035 ( .IN1(\ram[152][2] ), .IN2(n311), .IN3(n723), .IN4(datain[2]), 
        .Q(n2854) );
  AO22X1 U1036 ( .IN1(\ram[152][3] ), .IN2(n311), .IN3(n723), .IN4(datain[3]), 
        .Q(n2855) );
  AO22X1 U1037 ( .IN1(\ram[152][4] ), .IN2(n311), .IN3(n723), .IN4(datain[4]), 
        .Q(n2856) );
  AO22X1 U1038 ( .IN1(\ram[152][5] ), .IN2(n311), .IN3(n723), .IN4(datain[5]), 
        .Q(n2857) );
  AO22X1 U1039 ( .IN1(\ram[152][6] ), .IN2(n311), .IN3(n723), .IN4(datain[6]), 
        .Q(n2858) );
  AO22X1 U1040 ( .IN1(\ram[152][7] ), .IN2(n311), .IN3(n723), .IN4(datain[7]), 
        .Q(n2859) );
  AO22X1 U1043 ( .IN1(\ram[151][0] ), .IN2(n314), .IN3(n576), .IN4(datain[0]), 
        .Q(n2860) );
  AO22X1 U1044 ( .IN1(\ram[151][1] ), .IN2(n314), .IN3(n576), .IN4(datain[1]), 
        .Q(n2861) );
  AO22X1 U1045 ( .IN1(\ram[151][2] ), .IN2(n314), .IN3(n576), .IN4(datain[2]), 
        .Q(n2862) );
  AO22X1 U1046 ( .IN1(\ram[151][3] ), .IN2(n314), .IN3(n576), .IN4(datain[3]), 
        .Q(n2863) );
  AO22X1 U1047 ( .IN1(\ram[151][4] ), .IN2(n314), .IN3(n576), .IN4(datain[4]), 
        .Q(n2864) );
  AO22X1 U1048 ( .IN1(\ram[151][5] ), .IN2(n314), .IN3(n576), .IN4(datain[5]), 
        .Q(n2865) );
  AO22X1 U1049 ( .IN1(\ram[151][6] ), .IN2(n314), .IN3(n576), .IN4(datain[6]), 
        .Q(n2866) );
  AO22X1 U1050 ( .IN1(\ram[151][7] ), .IN2(n314), .IN3(n576), .IN4(datain[7]), 
        .Q(n2867) );
  AO22X1 U1053 ( .IN1(\ram[150][0] ), .IN2(n317), .IN3(n4163), .IN4(datain[0]), 
        .Q(n2868) );
  AO22X1 U1054 ( .IN1(\ram[150][1] ), .IN2(n317), .IN3(n4163), .IN4(datain[1]), 
        .Q(n2869) );
  AO22X1 U1055 ( .IN1(\ram[150][2] ), .IN2(n317), .IN3(n4163), .IN4(datain[2]), 
        .Q(n2870) );
  AO22X1 U1056 ( .IN1(\ram[150][3] ), .IN2(n317), .IN3(n4163), .IN4(datain[3]), 
        .Q(n2871) );
  AO22X1 U1057 ( .IN1(\ram[150][4] ), .IN2(n317), .IN3(n4163), .IN4(datain[4]), 
        .Q(n2872) );
  AO22X1 U1058 ( .IN1(\ram[150][5] ), .IN2(n317), .IN3(n4163), .IN4(datain[5]), 
        .Q(n2873) );
  AO22X1 U1059 ( .IN1(\ram[150][6] ), .IN2(n317), .IN3(n4163), .IN4(datain[6]), 
        .Q(n2874) );
  AO22X1 U1060 ( .IN1(\ram[150][7] ), .IN2(n317), .IN3(n4163), .IN4(datain[7]), 
        .Q(n2875) );
  AO22X1 U1063 ( .IN1(\ram[149][0] ), .IN2(n320), .IN3(n672), .IN4(datain[0]), 
        .Q(n2876) );
  AO22X1 U1064 ( .IN1(\ram[149][1] ), .IN2(n320), .IN3(n672), .IN4(datain[1]), 
        .Q(n2877) );
  AO22X1 U1065 ( .IN1(\ram[149][2] ), .IN2(n320), .IN3(n672), .IN4(datain[2]), 
        .Q(n2878) );
  AO22X1 U1066 ( .IN1(\ram[149][3] ), .IN2(n320), .IN3(n672), .IN4(datain[3]), 
        .Q(n2879) );
  AO22X1 U1067 ( .IN1(\ram[149][4] ), .IN2(n320), .IN3(n672), .IN4(datain[4]), 
        .Q(n2880) );
  AO22X1 U1068 ( .IN1(\ram[149][5] ), .IN2(n320), .IN3(n672), .IN4(datain[5]), 
        .Q(n2881) );
  AO22X1 U1069 ( .IN1(\ram[149][6] ), .IN2(n320), .IN3(n672), .IN4(datain[6]), 
        .Q(n2882) );
  AO22X1 U1070 ( .IN1(\ram[149][7] ), .IN2(n320), .IN3(n672), .IN4(datain[7]), 
        .Q(n2883) );
  AO22X1 U1073 ( .IN1(\ram[148][0] ), .IN2(n323), .IN3(n4115), .IN4(datain[0]), 
        .Q(n2884) );
  AO22X1 U1074 ( .IN1(\ram[148][1] ), .IN2(n323), .IN3(n4115), .IN4(datain[1]), 
        .Q(n2885) );
  AO22X1 U1075 ( .IN1(\ram[148][2] ), .IN2(n323), .IN3(n4115), .IN4(datain[2]), 
        .Q(n2886) );
  AO22X1 U1076 ( .IN1(\ram[148][3] ), .IN2(n323), .IN3(n4115), .IN4(datain[3]), 
        .Q(n2887) );
  AO22X1 U1077 ( .IN1(\ram[148][4] ), .IN2(n323), .IN3(n4115), .IN4(datain[4]), 
        .Q(n2888) );
  AO22X1 U1078 ( .IN1(\ram[148][5] ), .IN2(n323), .IN3(n4115), .IN4(datain[5]), 
        .Q(n2889) );
  AO22X1 U1079 ( .IN1(\ram[148][6] ), .IN2(n323), .IN3(n4115), .IN4(datain[6]), 
        .Q(n2890) );
  AO22X1 U1080 ( .IN1(\ram[148][7] ), .IN2(n323), .IN3(n4115), .IN4(datain[7]), 
        .Q(n2891) );
  AO22X1 U1083 ( .IN1(\ram[147][0] ), .IN2(n326), .IN3(n528), .IN4(datain[0]), 
        .Q(n2892) );
  AO22X1 U1084 ( .IN1(\ram[147][1] ), .IN2(n326), .IN3(n528), .IN4(datain[1]), 
        .Q(n2893) );
  AO22X1 U1085 ( .IN1(\ram[147][2] ), .IN2(n326), .IN3(n528), .IN4(datain[2]), 
        .Q(n2894) );
  AO22X1 U1086 ( .IN1(\ram[147][3] ), .IN2(n326), .IN3(n528), .IN4(datain[3]), 
        .Q(n2895) );
  AO22X1 U1087 ( .IN1(\ram[147][4] ), .IN2(n326), .IN3(n528), .IN4(datain[4]), 
        .Q(n2896) );
  AO22X1 U1088 ( .IN1(\ram[147][5] ), .IN2(n326), .IN3(n528), .IN4(datain[5]), 
        .Q(n2897) );
  AO22X1 U1089 ( .IN1(\ram[147][6] ), .IN2(n326), .IN3(n528), .IN4(datain[6]), 
        .Q(n2898) );
  AO22X1 U1090 ( .IN1(\ram[147][7] ), .IN2(n326), .IN3(n528), .IN4(datain[7]), 
        .Q(n2899) );
  AO22X1 U1093 ( .IN1(\ram[146][0] ), .IN2(n329), .IN3(n4147), .IN4(datain[0]), 
        .Q(n2900) );
  AO22X1 U1094 ( .IN1(\ram[146][1] ), .IN2(n329), .IN3(n4147), .IN4(datain[1]), 
        .Q(n2901) );
  AO22X1 U1095 ( .IN1(\ram[146][2] ), .IN2(n329), .IN3(n4147), .IN4(datain[2]), 
        .Q(n2902) );
  AO22X1 U1096 ( .IN1(\ram[146][3] ), .IN2(n329), .IN3(n4147), .IN4(datain[3]), 
        .Q(n2903) );
  AO22X1 U1097 ( .IN1(\ram[146][4] ), .IN2(n329), .IN3(n4147), .IN4(datain[4]), 
        .Q(n2904) );
  AO22X1 U1098 ( .IN1(\ram[146][5] ), .IN2(n329), .IN3(n4147), .IN4(datain[5]), 
        .Q(n2905) );
  AO22X1 U1099 ( .IN1(\ram[146][6] ), .IN2(n329), .IN3(n4147), .IN4(datain[6]), 
        .Q(n2906) );
  AO22X1 U1100 ( .IN1(\ram[146][7] ), .IN2(n329), .IN3(n4147), .IN4(datain[7]), 
        .Q(n2907) );
  AO22X1 U1103 ( .IN1(\ram[145][0] ), .IN2(n332), .IN3(n624), .IN4(datain[0]), 
        .Q(n2908) );
  AO22X1 U1104 ( .IN1(\ram[145][1] ), .IN2(n332), .IN3(n624), .IN4(datain[1]), 
        .Q(n2909) );
  AO22X1 U1105 ( .IN1(\ram[145][2] ), .IN2(n332), .IN3(n624), .IN4(datain[2]), 
        .Q(n2910) );
  AO22X1 U1106 ( .IN1(\ram[145][3] ), .IN2(n332), .IN3(n624), .IN4(datain[3]), 
        .Q(n2911) );
  AO22X1 U1107 ( .IN1(\ram[145][4] ), .IN2(n332), .IN3(n624), .IN4(datain[4]), 
        .Q(n2912) );
  AO22X1 U1108 ( .IN1(\ram[145][5] ), .IN2(n332), .IN3(n624), .IN4(datain[5]), 
        .Q(n2913) );
  AO22X1 U1109 ( .IN1(\ram[145][6] ), .IN2(n332), .IN3(n624), .IN4(datain[6]), 
        .Q(n2914) );
  AO22X1 U1110 ( .IN1(\ram[145][7] ), .IN2(n332), .IN3(n624), .IN4(datain[7]), 
        .Q(n2915) );
  AO22X1 U1113 ( .IN1(\ram[144][0] ), .IN2(n335), .IN3(n4130), .IN4(datain[0]), 
        .Q(n2916) );
  AO22X1 U1114 ( .IN1(\ram[144][1] ), .IN2(n335), .IN3(n4130), .IN4(datain[1]), 
        .Q(n2917) );
  AO22X1 U1115 ( .IN1(\ram[144][2] ), .IN2(n335), .IN3(n4130), .IN4(datain[2]), 
        .Q(n2918) );
  AO22X1 U1116 ( .IN1(\ram[144][3] ), .IN2(n335), .IN3(n4130), .IN4(datain[3]), 
        .Q(n2919) );
  AO22X1 U1117 ( .IN1(\ram[144][4] ), .IN2(n335), .IN3(n4130), .IN4(datain[4]), 
        .Q(n2920) );
  AO22X1 U1118 ( .IN1(\ram[144][5] ), .IN2(n335), .IN3(n4130), .IN4(datain[5]), 
        .Q(n2921) );
  AO22X1 U1119 ( .IN1(\ram[144][6] ), .IN2(n335), .IN3(n4130), .IN4(datain[6]), 
        .Q(n2922) );
  AO22X1 U1120 ( .IN1(\ram[144][7] ), .IN2(n335), .IN3(n4130), .IN4(datain[7]), 
        .Q(n2923) );
  AO22X1 U1123 ( .IN1(\ram[143][0] ), .IN2(n338), .IN3(n381), .IN4(datain[0]), 
        .Q(n2924) );
  AO22X1 U1124 ( .IN1(\ram[143][1] ), .IN2(n338), .IN3(n381), .IN4(datain[1]), 
        .Q(n2925) );
  AO22X1 U1125 ( .IN1(\ram[143][2] ), .IN2(n338), .IN3(n381), .IN4(datain[2]), 
        .Q(n2926) );
  AO22X1 U1126 ( .IN1(\ram[143][3] ), .IN2(n338), .IN3(n381), .IN4(datain[3]), 
        .Q(n2927) );
  AO22X1 U1127 ( .IN1(\ram[143][4] ), .IN2(n338), .IN3(n381), .IN4(datain[4]), 
        .Q(n2928) );
  AO22X1 U1128 ( .IN1(\ram[143][5] ), .IN2(n338), .IN3(n381), .IN4(datain[5]), 
        .Q(n2929) );
  AO22X1 U1129 ( .IN1(\ram[143][6] ), .IN2(n338), .IN3(n381), .IN4(datain[6]), 
        .Q(n2930) );
  AO22X1 U1130 ( .IN1(\ram[143][7] ), .IN2(n338), .IN3(n381), .IN4(datain[7]), 
        .Q(n2931) );
  AO22X1 U1133 ( .IN1(\ram[142][0] ), .IN2(n341), .IN3(n4101), .IN4(datain[0]), 
        .Q(n2932) );
  AO22X1 U1134 ( .IN1(\ram[142][1] ), .IN2(n341), .IN3(n4101), .IN4(datain[1]), 
        .Q(n2933) );
  AO22X1 U1135 ( .IN1(\ram[142][2] ), .IN2(n341), .IN3(n4101), .IN4(datain[2]), 
        .Q(n2934) );
  AO22X1 U1136 ( .IN1(\ram[142][3] ), .IN2(n341), .IN3(n4101), .IN4(datain[3]), 
        .Q(n2935) );
  AO22X1 U1137 ( .IN1(\ram[142][4] ), .IN2(n341), .IN3(n4101), .IN4(datain[4]), 
        .Q(n2936) );
  AO22X1 U1138 ( .IN1(\ram[142][5] ), .IN2(n341), .IN3(n4101), .IN4(datain[5]), 
        .Q(n2937) );
  AO22X1 U1139 ( .IN1(\ram[142][6] ), .IN2(n341), .IN3(n4101), .IN4(datain[6]), 
        .Q(n2938) );
  AO22X1 U1140 ( .IN1(\ram[142][7] ), .IN2(n341), .IN3(n4101), .IN4(datain[7]), 
        .Q(n2939) );
  AO22X1 U1143 ( .IN1(\ram[141][0] ), .IN2(n344), .IN3(n486), .IN4(datain[0]), 
        .Q(n2940) );
  AO22X1 U1144 ( .IN1(\ram[141][1] ), .IN2(n344), .IN3(n486), .IN4(datain[1]), 
        .Q(n2941) );
  AO22X1 U1145 ( .IN1(\ram[141][2] ), .IN2(n344), .IN3(n486), .IN4(datain[2]), 
        .Q(n2942) );
  AO22X1 U1146 ( .IN1(\ram[141][3] ), .IN2(n344), .IN3(n486), .IN4(datain[3]), 
        .Q(n2943) );
  AO22X1 U1147 ( .IN1(\ram[141][4] ), .IN2(n344), .IN3(n486), .IN4(datain[4]), 
        .Q(n2944) );
  AO22X1 U1148 ( .IN1(\ram[141][5] ), .IN2(n344), .IN3(n486), .IN4(datain[5]), 
        .Q(n2945) );
  AO22X1 U1149 ( .IN1(\ram[141][6] ), .IN2(n344), .IN3(n486), .IN4(datain[6]), 
        .Q(n2946) );
  AO22X1 U1150 ( .IN1(\ram[141][7] ), .IN2(n344), .IN3(n486), .IN4(datain[7]), 
        .Q(n2947) );
  AO22X1 U1153 ( .IN1(\ram[140][0] ), .IN2(n347), .IN3(n770), .IN4(datain[0]), 
        .Q(n2948) );
  AO22X1 U1154 ( .IN1(\ram[140][1] ), .IN2(n347), .IN3(n770), .IN4(datain[1]), 
        .Q(n2949) );
  AO22X1 U1155 ( .IN1(\ram[140][2] ), .IN2(n347), .IN3(n770), .IN4(datain[2]), 
        .Q(n2950) );
  AO22X1 U1156 ( .IN1(\ram[140][3] ), .IN2(n347), .IN3(n770), .IN4(datain[3]), 
        .Q(n2951) );
  AO22X1 U1157 ( .IN1(\ram[140][4] ), .IN2(n347), .IN3(n770), .IN4(datain[4]), 
        .Q(n2952) );
  AO22X1 U1158 ( .IN1(\ram[140][5] ), .IN2(n347), .IN3(n770), .IN4(datain[5]), 
        .Q(n2953) );
  AO22X1 U1159 ( .IN1(\ram[140][6] ), .IN2(n347), .IN3(n770), .IN4(datain[6]), 
        .Q(n2954) );
  AO22X1 U1160 ( .IN1(\ram[140][7] ), .IN2(n347), .IN3(n770), .IN4(datain[7]), 
        .Q(n2955) );
  AO22X1 U1163 ( .IN1(\ram[139][0] ), .IN2(n350), .IN3(n336), .IN4(datain[0]), 
        .Q(n2956) );
  AO22X1 U1164 ( .IN1(\ram[139][1] ), .IN2(n350), .IN3(n336), .IN4(datain[1]), 
        .Q(n2957) );
  AO22X1 U1165 ( .IN1(\ram[139][2] ), .IN2(n350), .IN3(n336), .IN4(datain[2]), 
        .Q(n2958) );
  AO22X1 U1166 ( .IN1(\ram[139][3] ), .IN2(n350), .IN3(n336), .IN4(datain[3]), 
        .Q(n2959) );
  AO22X1 U1167 ( .IN1(\ram[139][4] ), .IN2(n350), .IN3(n336), .IN4(datain[4]), 
        .Q(n2960) );
  AO22X1 U1168 ( .IN1(\ram[139][5] ), .IN2(n350), .IN3(n336), .IN4(datain[5]), 
        .Q(n2961) );
  AO22X1 U1169 ( .IN1(\ram[139][6] ), .IN2(n350), .IN3(n336), .IN4(datain[6]), 
        .Q(n2962) );
  AO22X1 U1170 ( .IN1(\ram[139][7] ), .IN2(n350), .IN3(n336), .IN4(datain[7]), 
        .Q(n2963) );
  AO22X1 U1173 ( .IN1(\ram[138][0] ), .IN2(n353), .IN3(n4084), .IN4(datain[0]), 
        .Q(n2964) );
  AO22X1 U1174 ( .IN1(\ram[138][1] ), .IN2(n353), .IN3(n4084), .IN4(datain[1]), 
        .Q(n2965) );
  AO22X1 U1175 ( .IN1(\ram[138][2] ), .IN2(n353), .IN3(n4084), .IN4(datain[2]), 
        .Q(n2966) );
  AO22X1 U1176 ( .IN1(\ram[138][3] ), .IN2(n353), .IN3(n4084), .IN4(datain[3]), 
        .Q(n2967) );
  AO22X1 U1177 ( .IN1(\ram[138][4] ), .IN2(n353), .IN3(n4084), .IN4(datain[4]), 
        .Q(n2968) );
  AO22X1 U1178 ( .IN1(\ram[138][5] ), .IN2(n353), .IN3(n4084), .IN4(datain[5]), 
        .Q(n2969) );
  AO22X1 U1179 ( .IN1(\ram[138][6] ), .IN2(n353), .IN3(n4084), .IN4(datain[6]), 
        .Q(n2970) );
  AO22X1 U1180 ( .IN1(\ram[138][7] ), .IN2(n353), .IN3(n4084), .IN4(datain[7]), 
        .Q(n2971) );
  AO22X1 U1183 ( .IN1(\ram[137][0] ), .IN2(n356), .IN3(n435), .IN4(datain[0]), 
        .Q(n2972) );
  AO22X1 U1184 ( .IN1(\ram[137][1] ), .IN2(n356), .IN3(n435), .IN4(datain[1]), 
        .Q(n2973) );
  AO22X1 U1185 ( .IN1(\ram[137][2] ), .IN2(n356), .IN3(n435), .IN4(datain[2]), 
        .Q(n2974) );
  AO22X1 U1186 ( .IN1(\ram[137][3] ), .IN2(n356), .IN3(n435), .IN4(datain[3]), 
        .Q(n2975) );
  AO22X1 U1187 ( .IN1(\ram[137][4] ), .IN2(n356), .IN3(n435), .IN4(datain[4]), 
        .Q(n2976) );
  AO22X1 U1188 ( .IN1(\ram[137][5] ), .IN2(n356), .IN3(n435), .IN4(datain[5]), 
        .Q(n2977) );
  AO22X1 U1189 ( .IN1(\ram[137][6] ), .IN2(n356), .IN3(n435), .IN4(datain[6]), 
        .Q(n2978) );
  AO22X1 U1190 ( .IN1(\ram[137][7] ), .IN2(n356), .IN3(n435), .IN4(datain[7]), 
        .Q(n2979) );
  AO22X1 U1193 ( .IN1(\ram[136][0] ), .IN2(n359), .IN3(n726), .IN4(datain[0]), 
        .Q(n2980) );
  AO22X1 U1194 ( .IN1(\ram[136][1] ), .IN2(n359), .IN3(n726), .IN4(datain[1]), 
        .Q(n2981) );
  AO22X1 U1195 ( .IN1(\ram[136][2] ), .IN2(n359), .IN3(n726), .IN4(datain[2]), 
        .Q(n2982) );
  AO22X1 U1196 ( .IN1(\ram[136][3] ), .IN2(n359), .IN3(n726), .IN4(datain[3]), 
        .Q(n2983) );
  AO22X1 U1197 ( .IN1(\ram[136][4] ), .IN2(n359), .IN3(n726), .IN4(datain[4]), 
        .Q(n2984) );
  AO22X1 U1198 ( .IN1(\ram[136][5] ), .IN2(n359), .IN3(n726), .IN4(datain[5]), 
        .Q(n2985) );
  AO22X1 U1199 ( .IN1(\ram[136][6] ), .IN2(n359), .IN3(n726), .IN4(datain[6]), 
        .Q(n2986) );
  AO22X1 U1200 ( .IN1(\ram[136][7] ), .IN2(n359), .IN3(n726), .IN4(datain[7]), 
        .Q(n2987) );
  AO22X1 U1203 ( .IN1(\ram[135][0] ), .IN2(n362), .IN3(n579), .IN4(datain[0]), 
        .Q(n2988) );
  AO22X1 U1204 ( .IN1(\ram[135][1] ), .IN2(n362), .IN3(n579), .IN4(datain[1]), 
        .Q(n2989) );
  AO22X1 U1205 ( .IN1(\ram[135][2] ), .IN2(n362), .IN3(n579), .IN4(datain[2]), 
        .Q(n2990) );
  AO22X1 U1206 ( .IN1(\ram[135][3] ), .IN2(n362), .IN3(n579), .IN4(datain[3]), 
        .Q(n2991) );
  AO22X1 U1207 ( .IN1(\ram[135][4] ), .IN2(n362), .IN3(n579), .IN4(datain[4]), 
        .Q(n2992) );
  AO22X1 U1208 ( .IN1(\ram[135][5] ), .IN2(n362), .IN3(n579), .IN4(datain[5]), 
        .Q(n2993) );
  AO22X1 U1209 ( .IN1(\ram[135][6] ), .IN2(n362), .IN3(n579), .IN4(datain[6]), 
        .Q(n2994) );
  AO22X1 U1210 ( .IN1(\ram[135][7] ), .IN2(n362), .IN3(n579), .IN4(datain[7]), 
        .Q(n2995) );
  AO22X1 U1213 ( .IN1(\ram[134][0] ), .IN2(n365), .IN3(n4164), .IN4(datain[0]), 
        .Q(n2996) );
  AO22X1 U1214 ( .IN1(\ram[134][1] ), .IN2(n365), .IN3(n4164), .IN4(datain[1]), 
        .Q(n2997) );
  AO22X1 U1215 ( .IN1(\ram[134][2] ), .IN2(n365), .IN3(n4164), .IN4(datain[2]), 
        .Q(n2998) );
  AO22X1 U1216 ( .IN1(\ram[134][3] ), .IN2(n365), .IN3(n4164), .IN4(datain[3]), 
        .Q(n2999) );
  AO22X1 U1217 ( .IN1(\ram[134][4] ), .IN2(n365), .IN3(n4164), .IN4(datain[4]), 
        .Q(n3000) );
  AO22X1 U1218 ( .IN1(\ram[134][5] ), .IN2(n365), .IN3(n4164), .IN4(datain[5]), 
        .Q(n3001) );
  AO22X1 U1219 ( .IN1(\ram[134][6] ), .IN2(n365), .IN3(n4164), .IN4(datain[6]), 
        .Q(n3002) );
  AO22X1 U1220 ( .IN1(\ram[134][7] ), .IN2(n365), .IN3(n4164), .IN4(datain[7]), 
        .Q(n3003) );
  AO22X1 U1223 ( .IN1(\ram[133][0] ), .IN2(n368), .IN3(n675), .IN4(datain[0]), 
        .Q(n3004) );
  AO22X1 U1224 ( .IN1(\ram[133][1] ), .IN2(n368), .IN3(n675), .IN4(datain[1]), 
        .Q(n3005) );
  AO22X1 U1225 ( .IN1(\ram[133][2] ), .IN2(n368), .IN3(n675), .IN4(datain[2]), 
        .Q(n3006) );
  AO22X1 U1226 ( .IN1(\ram[133][3] ), .IN2(n368), .IN3(n675), .IN4(datain[3]), 
        .Q(n3007) );
  AO22X1 U1227 ( .IN1(\ram[133][4] ), .IN2(n368), .IN3(n675), .IN4(datain[4]), 
        .Q(n3008) );
  AO22X1 U1228 ( .IN1(\ram[133][5] ), .IN2(n368), .IN3(n675), .IN4(datain[5]), 
        .Q(n3009) );
  AO22X1 U1229 ( .IN1(\ram[133][6] ), .IN2(n368), .IN3(n675), .IN4(datain[6]), 
        .Q(n3010) );
  AO22X1 U1230 ( .IN1(\ram[133][7] ), .IN2(n368), .IN3(n675), .IN4(datain[7]), 
        .Q(n3011) );
  AO22X1 U1233 ( .IN1(\ram[132][0] ), .IN2(n371), .IN3(n4116), .IN4(datain[0]), 
        .Q(n3012) );
  AO22X1 U1234 ( .IN1(\ram[132][1] ), .IN2(n371), .IN3(n4116), .IN4(datain[1]), 
        .Q(n3013) );
  AO22X1 U1235 ( .IN1(\ram[132][2] ), .IN2(n371), .IN3(n4116), .IN4(datain[2]), 
        .Q(n3014) );
  AO22X1 U1236 ( .IN1(\ram[132][3] ), .IN2(n371), .IN3(n4116), .IN4(datain[3]), 
        .Q(n3015) );
  AO22X1 U1237 ( .IN1(\ram[132][4] ), .IN2(n371), .IN3(n4116), .IN4(datain[4]), 
        .Q(n3016) );
  AO22X1 U1238 ( .IN1(\ram[132][5] ), .IN2(n371), .IN3(n4116), .IN4(datain[5]), 
        .Q(n3017) );
  AO22X1 U1239 ( .IN1(\ram[132][6] ), .IN2(n371), .IN3(n4116), .IN4(datain[6]), 
        .Q(n3018) );
  AO22X1 U1240 ( .IN1(\ram[132][7] ), .IN2(n371), .IN3(n4116), .IN4(datain[7]), 
        .Q(n3019) );
  AO22X1 U1243 ( .IN1(\ram[131][0] ), .IN2(n374), .IN3(n531), .IN4(n63), .Q(
        n3020) );
  AO22X1 U1244 ( .IN1(\ram[131][1] ), .IN2(n374), .IN3(n531), .IN4(n96), .Q(
        n3021) );
  AO22X1 U1245 ( .IN1(\ram[131][2] ), .IN2(n374), .IN3(n531), .IN4(n129), .Q(
        n3022) );
  AO22X1 U1246 ( .IN1(\ram[131][3] ), .IN2(n374), .IN3(n531), .IN4(n162), .Q(
        n3023) );
  AO22X1 U1247 ( .IN1(\ram[131][4] ), .IN2(n374), .IN3(n531), .IN4(n195), .Q(
        n3024) );
  AO22X1 U1248 ( .IN1(\ram[131][5] ), .IN2(n374), .IN3(n531), .IN4(n228), .Q(
        n3025) );
  AO22X1 U1249 ( .IN1(\ram[131][6] ), .IN2(n374), .IN3(n531), .IN4(n261), .Q(
        n3026) );
  AO22X1 U1250 ( .IN1(\ram[131][7] ), .IN2(n374), .IN3(n531), .IN4(n294), .Q(
        n3027) );
  AO22X1 U1253 ( .IN1(\ram[130][0] ), .IN2(n377), .IN3(n4148), .IN4(n63), .Q(
        n3028) );
  AO22X1 U1254 ( .IN1(\ram[130][1] ), .IN2(n377), .IN3(n4148), .IN4(n96), .Q(
        n3029) );
  AO22X1 U1255 ( .IN1(\ram[130][2] ), .IN2(n377), .IN3(n4148), .IN4(n129), .Q(
        n3030) );
  AO22X1 U1256 ( .IN1(\ram[130][3] ), .IN2(n377), .IN3(n4148), .IN4(n162), .Q(
        n3031) );
  AO22X1 U1257 ( .IN1(\ram[130][4] ), .IN2(n377), .IN3(n4148), .IN4(n195), .Q(
        n3032) );
  AO22X1 U1258 ( .IN1(\ram[130][5] ), .IN2(n377), .IN3(n4148), .IN4(n228), .Q(
        n3033) );
  AO22X1 U1259 ( .IN1(\ram[130][6] ), .IN2(n377), .IN3(n4148), .IN4(n261), .Q(
        n3034) );
  AO22X1 U1260 ( .IN1(\ram[130][7] ), .IN2(n377), .IN3(n4148), .IN4(n294), .Q(
        n3035) );
  AO22X1 U1263 ( .IN1(\ram[129][0] ), .IN2(n380), .IN3(n627), .IN4(n63), .Q(
        n3036) );
  AO22X1 U1264 ( .IN1(\ram[129][1] ), .IN2(n380), .IN3(n627), .IN4(n96), .Q(
        n3037) );
  AO22X1 U1265 ( .IN1(\ram[129][2] ), .IN2(n380), .IN3(n627), .IN4(n129), .Q(
        n3038) );
  AO22X1 U1266 ( .IN1(\ram[129][3] ), .IN2(n380), .IN3(n627), .IN4(n162), .Q(
        n3039) );
  AO22X1 U1267 ( .IN1(\ram[129][4] ), .IN2(n380), .IN3(n627), .IN4(n195), .Q(
        n3040) );
  AO22X1 U1268 ( .IN1(\ram[129][5] ), .IN2(n380), .IN3(n627), .IN4(n228), .Q(
        n3041) );
  AO22X1 U1269 ( .IN1(\ram[129][6] ), .IN2(n380), .IN3(n627), .IN4(n261), .Q(
        n3042) );
  AO22X1 U1270 ( .IN1(\ram[129][7] ), .IN2(n380), .IN3(n627), .IN4(n294), .Q(
        n3043) );
  AO22X1 U1273 ( .IN1(\ram[128][0] ), .IN2(n383), .IN3(n4121), .IN4(n63), .Q(
        n3044) );
  AO22X1 U1274 ( .IN1(\ram[128][1] ), .IN2(n383), .IN3(n4121), .IN4(n96), .Q(
        n3045) );
  AO22X1 U1275 ( .IN1(\ram[128][2] ), .IN2(n383), .IN3(n4121), .IN4(n129), .Q(
        n3046) );
  AO22X1 U1276 ( .IN1(\ram[128][3] ), .IN2(n383), .IN3(n4121), .IN4(n162), .Q(
        n3047) );
  AO22X1 U1277 ( .IN1(\ram[128][4] ), .IN2(n383), .IN3(n4121), .IN4(n195), .Q(
        n3048) );
  AO22X1 U1278 ( .IN1(\ram[128][5] ), .IN2(n383), .IN3(n4121), .IN4(n228), .Q(
        n3049) );
  AO22X1 U1279 ( .IN1(\ram[128][6] ), .IN2(n383), .IN3(n4121), .IN4(n261), .Q(
        n3050) );
  AO22X1 U1280 ( .IN1(\ram[128][7] ), .IN2(n383), .IN3(n4121), .IN4(n294), .Q(
        n3051) );
  AO22X1 U1283 ( .IN1(\ram[127][0] ), .IN2(n386), .IN3(n354), .IN4(n63), .Q(
        n3052) );
  AO22X1 U1284 ( .IN1(\ram[127][1] ), .IN2(n386), .IN3(n354), .IN4(n96), .Q(
        n3053) );
  AO22X1 U1285 ( .IN1(\ram[127][2] ), .IN2(n386), .IN3(n354), .IN4(n129), .Q(
        n3054) );
  AO22X1 U1286 ( .IN1(\ram[127][3] ), .IN2(n386), .IN3(n354), .IN4(n162), .Q(
        n3055) );
  AO22X1 U1287 ( .IN1(\ram[127][4] ), .IN2(n386), .IN3(n354), .IN4(n195), .Q(
        n3056) );
  AO22X1 U1288 ( .IN1(\ram[127][5] ), .IN2(n386), .IN3(n354), .IN4(n228), .Q(
        n3057) );
  AO22X1 U1289 ( .IN1(\ram[127][6] ), .IN2(n386), .IN3(n354), .IN4(n261), .Q(
        n3058) );
  AO22X1 U1290 ( .IN1(\ram[127][7] ), .IN2(n386), .IN3(n354), .IN4(n294), .Q(
        n3059) );
  AO22X1 U1293 ( .IN1(\ram[126][0] ), .IN2(n389), .IN3(n4092), .IN4(n63), .Q(
        n3060) );
  AO22X1 U1294 ( .IN1(\ram[126][1] ), .IN2(n389), .IN3(n4092), .IN4(n96), .Q(
        n3061) );
  AO22X1 U1295 ( .IN1(\ram[126][2] ), .IN2(n389), .IN3(n4092), .IN4(n129), .Q(
        n3062) );
  AO22X1 U1296 ( .IN1(\ram[126][3] ), .IN2(n389), .IN3(n4092), .IN4(n162), .Q(
        n3063) );
  AO22X1 U1297 ( .IN1(\ram[126][4] ), .IN2(n389), .IN3(n4092), .IN4(n195), .Q(
        n3064) );
  AO22X1 U1298 ( .IN1(\ram[126][5] ), .IN2(n389), .IN3(n4092), .IN4(n228), .Q(
        n3065) );
  AO22X1 U1299 ( .IN1(\ram[126][6] ), .IN2(n389), .IN3(n4092), .IN4(n261), .Q(
        n3066) );
  AO22X1 U1300 ( .IN1(\ram[126][7] ), .IN2(n389), .IN3(n4092), .IN4(n294), .Q(
        n3067) );
  AO22X1 U1303 ( .IN1(\ram[125][0] ), .IN2(n392), .IN3(n459), .IN4(n63), .Q(
        n3068) );
  AO22X1 U1304 ( .IN1(\ram[125][1] ), .IN2(n392), .IN3(n459), .IN4(n96), .Q(
        n3069) );
  AO22X1 U1305 ( .IN1(\ram[125][2] ), .IN2(n392), .IN3(n459), .IN4(n129), .Q(
        n3070) );
  AO22X1 U1306 ( .IN1(\ram[125][3] ), .IN2(n392), .IN3(n459), .IN4(n162), .Q(
        n3071) );
  AO22X1 U1307 ( .IN1(\ram[125][4] ), .IN2(n392), .IN3(n459), .IN4(n195), .Q(
        n3072) );
  AO22X1 U1308 ( .IN1(\ram[125][5] ), .IN2(n392), .IN3(n459), .IN4(n228), .Q(
        n3073) );
  AO22X1 U1309 ( .IN1(\ram[125][6] ), .IN2(n392), .IN3(n459), .IN4(n261), .Q(
        n3074) );
  AO22X1 U1310 ( .IN1(\ram[125][7] ), .IN2(n392), .IN3(n459), .IN4(n294), .Q(
        n3075) );
  AO22X1 U1313 ( .IN1(\ram[124][0] ), .IN2(n395), .IN3(n741), .IN4(n63), .Q(
        n3076) );
  AO22X1 U1314 ( .IN1(\ram[124][1] ), .IN2(n395), .IN3(n741), .IN4(n96), .Q(
        n3077) );
  AO22X1 U1315 ( .IN1(\ram[124][2] ), .IN2(n395), .IN3(n741), .IN4(n129), .Q(
        n3078) );
  AO22X1 U1316 ( .IN1(\ram[124][3] ), .IN2(n395), .IN3(n741), .IN4(n162), .Q(
        n3079) );
  AO22X1 U1317 ( .IN1(\ram[124][4] ), .IN2(n395), .IN3(n741), .IN4(n195), .Q(
        n3080) );
  AO22X1 U1318 ( .IN1(\ram[124][5] ), .IN2(n395), .IN3(n741), .IN4(n228), .Q(
        n3081) );
  AO22X1 U1319 ( .IN1(\ram[124][6] ), .IN2(n395), .IN3(n741), .IN4(n261), .Q(
        n3082) );
  AO22X1 U1320 ( .IN1(\ram[124][7] ), .IN2(n395), .IN3(n741), .IN4(n294), .Q(
        n3083) );
  AO22X1 U1323 ( .IN1(\ram[123][0] ), .IN2(n398), .IN3(n306), .IN4(n63), .Q(
        n3084) );
  AO22X1 U1324 ( .IN1(\ram[123][1] ), .IN2(n398), .IN3(n306), .IN4(n96), .Q(
        n3085) );
  AO22X1 U1325 ( .IN1(\ram[123][2] ), .IN2(n398), .IN3(n306), .IN4(n129), .Q(
        n3086) );
  AO22X1 U1326 ( .IN1(\ram[123][3] ), .IN2(n398), .IN3(n306), .IN4(n162), .Q(
        n3087) );
  AO22X1 U1327 ( .IN1(\ram[123][4] ), .IN2(n398), .IN3(n306), .IN4(n195), .Q(
        n3088) );
  AO22X1 U1328 ( .IN1(\ram[123][5] ), .IN2(n398), .IN3(n306), .IN4(n228), .Q(
        n3089) );
  AO22X1 U1329 ( .IN1(\ram[123][6] ), .IN2(n398), .IN3(n306), .IN4(n261), .Q(
        n3090) );
  AO22X1 U1330 ( .IN1(\ram[123][7] ), .IN2(n398), .IN3(n306), .IN4(n294), .Q(
        n3091) );
  AO22X1 U1333 ( .IN1(\ram[122][0] ), .IN2(n401), .IN3(n2018), .IN4(n63), .Q(
        n3092) );
  AO22X1 U1334 ( .IN1(\ram[122][1] ), .IN2(n401), .IN3(n2018), .IN4(n96), .Q(
        n3093) );
  AO22X1 U1335 ( .IN1(\ram[122][2] ), .IN2(n401), .IN3(n2018), .IN4(n129), .Q(
        n3094) );
  AO22X1 U1336 ( .IN1(\ram[122][3] ), .IN2(n401), .IN3(n2018), .IN4(n162), .Q(
        n3095) );
  AO22X1 U1337 ( .IN1(\ram[122][4] ), .IN2(n401), .IN3(n2018), .IN4(n195), .Q(
        n3096) );
  AO22X1 U1338 ( .IN1(\ram[122][5] ), .IN2(n401), .IN3(n2018), .IN4(n228), .Q(
        n3097) );
  AO22X1 U1339 ( .IN1(\ram[122][6] ), .IN2(n401), .IN3(n2018), .IN4(n261), .Q(
        n3098) );
  AO22X1 U1340 ( .IN1(\ram[122][7] ), .IN2(n401), .IN3(n2018), .IN4(n294), .Q(
        n3099) );
  AO22X1 U1343 ( .IN1(\ram[121][0] ), .IN2(n404), .IN3(n405), .IN4(n63), .Q(
        n3100) );
  AO22X1 U1344 ( .IN1(\ram[121][1] ), .IN2(n404), .IN3(n405), .IN4(n96), .Q(
        n3101) );
  AO22X1 U1345 ( .IN1(\ram[121][2] ), .IN2(n404), .IN3(n405), .IN4(n129), .Q(
        n3102) );
  AO22X1 U1346 ( .IN1(\ram[121][3] ), .IN2(n404), .IN3(n405), .IN4(n162), .Q(
        n3103) );
  AO22X1 U1347 ( .IN1(\ram[121][4] ), .IN2(n404), .IN3(n405), .IN4(n195), .Q(
        n3104) );
  AO22X1 U1348 ( .IN1(\ram[121][5] ), .IN2(n404), .IN3(n405), .IN4(n228), .Q(
        n3105) );
  AO22X1 U1349 ( .IN1(\ram[121][6] ), .IN2(n404), .IN3(n405), .IN4(n261), .Q(
        n3106) );
  AO22X1 U1350 ( .IN1(\ram[121][7] ), .IN2(n404), .IN3(n405), .IN4(n294), .Q(
        n3107) );
  AO22X1 U1353 ( .IN1(\ram[120][0] ), .IN2(n407), .IN3(n693), .IN4(n63), .Q(
        n3108) );
  AO22X1 U1354 ( .IN1(\ram[120][1] ), .IN2(n407), .IN3(n693), .IN4(n96), .Q(
        n3109) );
  AO22X1 U1355 ( .IN1(\ram[120][2] ), .IN2(n407), .IN3(n693), .IN4(n129), .Q(
        n3110) );
  AO22X1 U1356 ( .IN1(\ram[120][3] ), .IN2(n407), .IN3(n693), .IN4(n162), .Q(
        n3111) );
  AO22X1 U1357 ( .IN1(\ram[120][4] ), .IN2(n407), .IN3(n693), .IN4(n195), .Q(
        n3112) );
  AO22X1 U1358 ( .IN1(\ram[120][5] ), .IN2(n407), .IN3(n693), .IN4(n228), .Q(
        n3113) );
  AO22X1 U1359 ( .IN1(\ram[120][6] ), .IN2(n407), .IN3(n693), .IN4(n261), .Q(
        n3114) );
  AO22X1 U1360 ( .IN1(\ram[120][7] ), .IN2(n407), .IN3(n693), .IN4(n294), .Q(
        n3115) );
  AO22X1 U1363 ( .IN1(\ram[119][0] ), .IN2(n410), .IN3(n546), .IN4(n60), .Q(
        n3116) );
  AO22X1 U1364 ( .IN1(\ram[119][1] ), .IN2(n410), .IN3(n546), .IN4(n93), .Q(
        n3117) );
  AO22X1 U1365 ( .IN1(\ram[119][2] ), .IN2(n410), .IN3(n546), .IN4(n126), .Q(
        n3118) );
  AO22X1 U1366 ( .IN1(\ram[119][3] ), .IN2(n410), .IN3(n546), .IN4(n159), .Q(
        n3119) );
  AO22X1 U1367 ( .IN1(\ram[119][4] ), .IN2(n410), .IN3(n546), .IN4(n192), .Q(
        n3120) );
  AO22X1 U1368 ( .IN1(\ram[119][5] ), .IN2(n410), .IN3(n546), .IN4(n225), .Q(
        n3121) );
  AO22X1 U1369 ( .IN1(\ram[119][6] ), .IN2(n410), .IN3(n546), .IN4(n258), .Q(
        n3122) );
  AO22X1 U1370 ( .IN1(\ram[119][7] ), .IN2(n410), .IN3(n546), .IN4(n291), .Q(
        n3123) );
  AO22X1 U1373 ( .IN1(\ram[118][0] ), .IN2(n413), .IN3(n4153), .IN4(n60), .Q(
        n3124) );
  AO22X1 U1374 ( .IN1(\ram[118][1] ), .IN2(n413), .IN3(n4153), .IN4(n93), .Q(
        n3125) );
  AO22X1 U1375 ( .IN1(\ram[118][2] ), .IN2(n413), .IN3(n4153), .IN4(n126), .Q(
        n3126) );
  AO22X1 U1376 ( .IN1(\ram[118][3] ), .IN2(n413), .IN3(n4153), .IN4(n159), .Q(
        n3127) );
  AO22X1 U1377 ( .IN1(\ram[118][4] ), .IN2(n413), .IN3(n4153), .IN4(n192), .Q(
        n3128) );
  AO22X1 U1378 ( .IN1(\ram[118][5] ), .IN2(n413), .IN3(n4153), .IN4(n225), .Q(
        n3129) );
  AO22X1 U1379 ( .IN1(\ram[118][6] ), .IN2(n413), .IN3(n4153), .IN4(n258), .Q(
        n3130) );
  AO22X1 U1380 ( .IN1(\ram[118][7] ), .IN2(n413), .IN3(n4153), .IN4(n291), .Q(
        n3131) );
  AO22X1 U1383 ( .IN1(\ram[117][0] ), .IN2(n416), .IN3(n642), .IN4(n60), .Q(
        n3132) );
  AO22X1 U1384 ( .IN1(\ram[117][1] ), .IN2(n416), .IN3(n642), .IN4(n93), .Q(
        n3133) );
  AO22X1 U1385 ( .IN1(\ram[117][2] ), .IN2(n416), .IN3(n642), .IN4(n126), .Q(
        n3134) );
  AO22X1 U1386 ( .IN1(\ram[117][3] ), .IN2(n416), .IN3(n642), .IN4(n159), .Q(
        n3135) );
  AO22X1 U1387 ( .IN1(\ram[117][4] ), .IN2(n416), .IN3(n642), .IN4(n192), .Q(
        n3136) );
  AO22X1 U1388 ( .IN1(\ram[117][5] ), .IN2(n416), .IN3(n642), .IN4(n225), .Q(
        n3137) );
  AO22X1 U1389 ( .IN1(\ram[117][6] ), .IN2(n416), .IN3(n642), .IN4(n258), .Q(
        n3138) );
  AO22X1 U1390 ( .IN1(\ram[117][7] ), .IN2(n416), .IN3(n642), .IN4(n291), .Q(
        n3139) );
  AO22X1 U1393 ( .IN1(\ram[116][0] ), .IN2(n419), .IN3(n4105), .IN4(n60), .Q(
        n3140) );
  AO22X1 U1394 ( .IN1(\ram[116][1] ), .IN2(n419), .IN3(n4105), .IN4(n93), .Q(
        n3141) );
  AO22X1 U1395 ( .IN1(\ram[116][2] ), .IN2(n419), .IN3(n4105), .IN4(n126), .Q(
        n3142) );
  AO22X1 U1396 ( .IN1(\ram[116][3] ), .IN2(n419), .IN3(n4105), .IN4(n159), .Q(
        n3143) );
  AO22X1 U1397 ( .IN1(\ram[116][4] ), .IN2(n419), .IN3(n4105), .IN4(n192), .Q(
        n3144) );
  AO22X1 U1398 ( .IN1(\ram[116][5] ), .IN2(n419), .IN3(n4105), .IN4(n225), .Q(
        n3145) );
  AO22X1 U1399 ( .IN1(\ram[116][6] ), .IN2(n419), .IN3(n4105), .IN4(n258), .Q(
        n3146) );
  AO22X1 U1400 ( .IN1(\ram[116][7] ), .IN2(n419), .IN3(n4105), .IN4(n291), .Q(
        n3147) );
  AO22X1 U1403 ( .IN1(\ram[115][0] ), .IN2(n422), .IN3(n498), .IN4(n60), .Q(
        n3148) );
  AO22X1 U1404 ( .IN1(\ram[115][1] ), .IN2(n422), .IN3(n498), .IN4(n93), .Q(
        n3149) );
  AO22X1 U1405 ( .IN1(\ram[115][2] ), .IN2(n422), .IN3(n498), .IN4(n126), .Q(
        n3150) );
  AO22X1 U1406 ( .IN1(\ram[115][3] ), .IN2(n422), .IN3(n498), .IN4(n159), .Q(
        n3151) );
  AO22X1 U1407 ( .IN1(\ram[115][4] ), .IN2(n422), .IN3(n498), .IN4(n192), .Q(
        n3152) );
  AO22X1 U1408 ( .IN1(\ram[115][5] ), .IN2(n422), .IN3(n498), .IN4(n225), .Q(
        n3153) );
  AO22X1 U1409 ( .IN1(\ram[115][6] ), .IN2(n422), .IN3(n498), .IN4(n258), .Q(
        n3154) );
  AO22X1 U1410 ( .IN1(\ram[115][7] ), .IN2(n422), .IN3(n498), .IN4(n291), .Q(
        n3155) );
  AO22X1 U1413 ( .IN1(\ram[114][0] ), .IN2(n425), .IN3(n4137), .IN4(n60), .Q(
        n3156) );
  AO22X1 U1414 ( .IN1(\ram[114][1] ), .IN2(n425), .IN3(n4137), .IN4(n93), .Q(
        n3157) );
  AO22X1 U1415 ( .IN1(\ram[114][2] ), .IN2(n425), .IN3(n4137), .IN4(n126), .Q(
        n3158) );
  AO22X1 U1416 ( .IN1(\ram[114][3] ), .IN2(n425), .IN3(n4137), .IN4(n159), .Q(
        n3159) );
  AO22X1 U1417 ( .IN1(\ram[114][4] ), .IN2(n425), .IN3(n4137), .IN4(n192), .Q(
        n3160) );
  AO22X1 U1418 ( .IN1(\ram[114][5] ), .IN2(n425), .IN3(n4137), .IN4(n225), .Q(
        n3161) );
  AO22X1 U1419 ( .IN1(\ram[114][6] ), .IN2(n425), .IN3(n4137), .IN4(n258), .Q(
        n3162) );
  AO22X1 U1420 ( .IN1(\ram[114][7] ), .IN2(n425), .IN3(n4137), .IN4(n291), .Q(
        n3163) );
  AO22X1 U1423 ( .IN1(\ram[113][0] ), .IN2(n428), .IN3(n594), .IN4(n60), .Q(
        n3164) );
  AO22X1 U1424 ( .IN1(\ram[113][1] ), .IN2(n428), .IN3(n594), .IN4(n93), .Q(
        n3165) );
  AO22X1 U1425 ( .IN1(\ram[113][2] ), .IN2(n428), .IN3(n594), .IN4(n126), .Q(
        n3166) );
  AO22X1 U1426 ( .IN1(\ram[113][3] ), .IN2(n428), .IN3(n594), .IN4(n159), .Q(
        n3167) );
  AO22X1 U1427 ( .IN1(\ram[113][4] ), .IN2(n428), .IN3(n594), .IN4(n192), .Q(
        n3168) );
  AO22X1 U1428 ( .IN1(\ram[113][5] ), .IN2(n428), .IN3(n594), .IN4(n225), .Q(
        n3169) );
  AO22X1 U1429 ( .IN1(\ram[113][6] ), .IN2(n428), .IN3(n594), .IN4(n258), .Q(
        n3170) );
  AO22X1 U1430 ( .IN1(\ram[113][7] ), .IN2(n428), .IN3(n594), .IN4(n291), .Q(
        n3171) );
  AO22X1 U1433 ( .IN1(\ram[112][0] ), .IN2(n431), .IN3(n4122), .IN4(n60), .Q(
        n3172) );
  AO22X1 U1434 ( .IN1(\ram[112][1] ), .IN2(n431), .IN3(n4122), .IN4(n93), .Q(
        n3173) );
  AO22X1 U1435 ( .IN1(\ram[112][2] ), .IN2(n431), .IN3(n4122), .IN4(n126), .Q(
        n3174) );
  AO22X1 U1436 ( .IN1(\ram[112][3] ), .IN2(n431), .IN3(n4122), .IN4(n159), .Q(
        n3175) );
  AO22X1 U1437 ( .IN1(\ram[112][4] ), .IN2(n431), .IN3(n4122), .IN4(n192), .Q(
        n3176) );
  AO22X1 U1438 ( .IN1(\ram[112][5] ), .IN2(n431), .IN3(n4122), .IN4(n225), .Q(
        n3177) );
  AO22X1 U1439 ( .IN1(\ram[112][6] ), .IN2(n431), .IN3(n4122), .IN4(n258), .Q(
        n3178) );
  AO22X1 U1440 ( .IN1(\ram[112][7] ), .IN2(n431), .IN3(n4122), .IN4(n291), .Q(
        n3179) );
  AO22X1 U1443 ( .IN1(\ram[111][0] ), .IN2(n434), .IN3(n357), .IN4(n60), .Q(
        n3180) );
  AO22X1 U1444 ( .IN1(\ram[111][1] ), .IN2(n434), .IN3(n357), .IN4(n93), .Q(
        n3181) );
  AO22X1 U1445 ( .IN1(\ram[111][2] ), .IN2(n434), .IN3(n357), .IN4(n126), .Q(
        n3182) );
  AO22X1 U1446 ( .IN1(\ram[111][3] ), .IN2(n434), .IN3(n357), .IN4(n159), .Q(
        n3183) );
  AO22X1 U1447 ( .IN1(\ram[111][4] ), .IN2(n434), .IN3(n357), .IN4(n192), .Q(
        n3184) );
  AO22X1 U1448 ( .IN1(\ram[111][5] ), .IN2(n434), .IN3(n357), .IN4(n225), .Q(
        n3185) );
  AO22X1 U1449 ( .IN1(\ram[111][6] ), .IN2(n434), .IN3(n357), .IN4(n258), .Q(
        n3186) );
  AO22X1 U1450 ( .IN1(\ram[111][7] ), .IN2(n434), .IN3(n357), .IN4(n291), .Q(
        n3187) );
  AO22X1 U1453 ( .IN1(\ram[110][0] ), .IN2(n437), .IN3(n4093), .IN4(n60), .Q(
        n3188) );
  AO22X1 U1454 ( .IN1(\ram[110][1] ), .IN2(n437), .IN3(n4093), .IN4(n93), .Q(
        n3189) );
  AO22X1 U1455 ( .IN1(\ram[110][2] ), .IN2(n437), .IN3(n4093), .IN4(n126), .Q(
        n3190) );
  AO22X1 U1456 ( .IN1(\ram[110][3] ), .IN2(n437), .IN3(n4093), .IN4(n159), .Q(
        n3191) );
  AO22X1 U1457 ( .IN1(\ram[110][4] ), .IN2(n437), .IN3(n4093), .IN4(n192), .Q(
        n3192) );
  AO22X1 U1458 ( .IN1(\ram[110][5] ), .IN2(n437), .IN3(n4093), .IN4(n225), .Q(
        n3193) );
  AO22X1 U1459 ( .IN1(\ram[110][6] ), .IN2(n437), .IN3(n4093), .IN4(n258), .Q(
        n3194) );
  AO22X1 U1460 ( .IN1(\ram[110][7] ), .IN2(n437), .IN3(n4093), .IN4(n291), .Q(
        n3195) );
  AO22X1 U1463 ( .IN1(\ram[109][0] ), .IN2(n440), .IN3(n462), .IN4(n60), .Q(
        n3196) );
  AO22X1 U1464 ( .IN1(\ram[109][1] ), .IN2(n440), .IN3(n462), .IN4(n93), .Q(
        n3197) );
  AO22X1 U1465 ( .IN1(\ram[109][2] ), .IN2(n440), .IN3(n462), .IN4(n126), .Q(
        n3198) );
  AO22X1 U1466 ( .IN1(\ram[109][3] ), .IN2(n440), .IN3(n462), .IN4(n159), .Q(
        n3199) );
  AO22X1 U1467 ( .IN1(\ram[109][4] ), .IN2(n440), .IN3(n462), .IN4(n192), .Q(
        n3200) );
  AO22X1 U1468 ( .IN1(\ram[109][5] ), .IN2(n440), .IN3(n462), .IN4(n225), .Q(
        n3201) );
  AO22X1 U1469 ( .IN1(\ram[109][6] ), .IN2(n440), .IN3(n462), .IN4(n258), .Q(
        n3202) );
  AO22X1 U1470 ( .IN1(\ram[109][7] ), .IN2(n440), .IN3(n462), .IN4(n291), .Q(
        n3203) );
  AO22X1 U1473 ( .IN1(\ram[108][0] ), .IN2(n443), .IN3(n744), .IN4(n60), .Q(
        n3204) );
  AO22X1 U1474 ( .IN1(\ram[108][1] ), .IN2(n443), .IN3(n744), .IN4(n93), .Q(
        n3205) );
  AO22X1 U1475 ( .IN1(\ram[108][2] ), .IN2(n443), .IN3(n744), .IN4(n126), .Q(
        n3206) );
  AO22X1 U1476 ( .IN1(\ram[108][3] ), .IN2(n443), .IN3(n744), .IN4(n159), .Q(
        n3207) );
  AO22X1 U1477 ( .IN1(\ram[108][4] ), .IN2(n443), .IN3(n744), .IN4(n192), .Q(
        n3208) );
  AO22X1 U1478 ( .IN1(\ram[108][5] ), .IN2(n443), .IN3(n744), .IN4(n225), .Q(
        n3209) );
  AO22X1 U1479 ( .IN1(\ram[108][6] ), .IN2(n443), .IN3(n744), .IN4(n258), .Q(
        n3210) );
  AO22X1 U1480 ( .IN1(\ram[108][7] ), .IN2(n443), .IN3(n744), .IN4(n291), .Q(
        n3211) );
  AO22X1 U1483 ( .IN1(\ram[107][0] ), .IN2(n446), .IN3(n309), .IN4(n57), .Q(
        n3212) );
  AO22X1 U1484 ( .IN1(\ram[107][1] ), .IN2(n446), .IN3(n309), .IN4(n90), .Q(
        n3213) );
  AO22X1 U1485 ( .IN1(\ram[107][2] ), .IN2(n446), .IN3(n309), .IN4(n123), .Q(
        n3214) );
  AO22X1 U1486 ( .IN1(\ram[107][3] ), .IN2(n446), .IN3(n309), .IN4(n156), .Q(
        n3215) );
  AO22X1 U1487 ( .IN1(\ram[107][4] ), .IN2(n446), .IN3(n309), .IN4(n189), .Q(
        n3216) );
  AO22X1 U1488 ( .IN1(\ram[107][5] ), .IN2(n446), .IN3(n309), .IN4(n222), .Q(
        n3217) );
  AO22X1 U1489 ( .IN1(\ram[107][6] ), .IN2(n446), .IN3(n309), .IN4(n255), .Q(
        n3218) );
  AO22X1 U1490 ( .IN1(\ram[107][7] ), .IN2(n446), .IN3(n309), .IN4(n288), .Q(
        n3219) );
  AO22X1 U1493 ( .IN1(\ram[106][0] ), .IN2(n449), .IN3(n2019), .IN4(n57), .Q(
        n3220) );
  AO22X1 U1494 ( .IN1(\ram[106][1] ), .IN2(n449), .IN3(n2019), .IN4(n90), .Q(
        n3221) );
  AO22X1 U1495 ( .IN1(\ram[106][2] ), .IN2(n449), .IN3(n2019), .IN4(n123), .Q(
        n3222) );
  AO22X1 U1496 ( .IN1(\ram[106][3] ), .IN2(n449), .IN3(n2019), .IN4(n156), .Q(
        n3223) );
  AO22X1 U1497 ( .IN1(\ram[106][4] ), .IN2(n449), .IN3(n2019), .IN4(n189), .Q(
        n3224) );
  AO22X1 U1498 ( .IN1(\ram[106][5] ), .IN2(n449), .IN3(n2019), .IN4(n222), .Q(
        n3225) );
  AO22X1 U1499 ( .IN1(\ram[106][6] ), .IN2(n449), .IN3(n2019), .IN4(n255), .Q(
        n3226) );
  AO22X1 U1500 ( .IN1(\ram[106][7] ), .IN2(n449), .IN3(n2019), .IN4(n288), .Q(
        n3227) );
  AO22X1 U1503 ( .IN1(\ram[105][0] ), .IN2(n452), .IN3(n408), .IN4(n57), .Q(
        n3228) );
  AO22X1 U1504 ( .IN1(\ram[105][1] ), .IN2(n452), .IN3(n408), .IN4(n90), .Q(
        n3229) );
  AO22X1 U1505 ( .IN1(\ram[105][2] ), .IN2(n452), .IN3(n408), .IN4(n123), .Q(
        n3230) );
  AO22X1 U1506 ( .IN1(\ram[105][3] ), .IN2(n452), .IN3(n408), .IN4(n156), .Q(
        n3231) );
  AO22X1 U1507 ( .IN1(\ram[105][4] ), .IN2(n452), .IN3(n408), .IN4(n189), .Q(
        n3232) );
  AO22X1 U1508 ( .IN1(\ram[105][5] ), .IN2(n452), .IN3(n408), .IN4(n222), .Q(
        n3233) );
  AO22X1 U1509 ( .IN1(\ram[105][6] ), .IN2(n452), .IN3(n408), .IN4(n255), .Q(
        n3234) );
  AO22X1 U1510 ( .IN1(\ram[105][7] ), .IN2(n452), .IN3(n408), .IN4(n288), .Q(
        n3235) );
  AO22X1 U1513 ( .IN1(\ram[104][0] ), .IN2(n455), .IN3(n696), .IN4(n57), .Q(
        n3236) );
  AO22X1 U1514 ( .IN1(\ram[104][1] ), .IN2(n455), .IN3(n696), .IN4(n90), .Q(
        n3237) );
  AO22X1 U1515 ( .IN1(\ram[104][2] ), .IN2(n455), .IN3(n696), .IN4(n123), .Q(
        n3238) );
  AO22X1 U1516 ( .IN1(\ram[104][3] ), .IN2(n455), .IN3(n696), .IN4(n156), .Q(
        n3239) );
  AO22X1 U1517 ( .IN1(\ram[104][4] ), .IN2(n455), .IN3(n696), .IN4(n189), .Q(
        n3240) );
  AO22X1 U1518 ( .IN1(\ram[104][5] ), .IN2(n455), .IN3(n696), .IN4(n222), .Q(
        n3241) );
  AO22X1 U1519 ( .IN1(\ram[104][6] ), .IN2(n455), .IN3(n696), .IN4(n255), .Q(
        n3242) );
  AO22X1 U1520 ( .IN1(\ram[104][7] ), .IN2(n455), .IN3(n696), .IN4(n288), .Q(
        n3243) );
  AO22X1 U1523 ( .IN1(\ram[103][0] ), .IN2(n458), .IN3(n549), .IN4(n57), .Q(
        n3244) );
  AO22X1 U1524 ( .IN1(\ram[103][1] ), .IN2(n458), .IN3(n549), .IN4(n90), .Q(
        n3245) );
  AO22X1 U1525 ( .IN1(\ram[103][2] ), .IN2(n458), .IN3(n549), .IN4(n123), .Q(
        n3246) );
  AO22X1 U1526 ( .IN1(\ram[103][3] ), .IN2(n458), .IN3(n549), .IN4(n156), .Q(
        n3247) );
  AO22X1 U1527 ( .IN1(\ram[103][4] ), .IN2(n458), .IN3(n549), .IN4(n189), .Q(
        n3248) );
  AO22X1 U1528 ( .IN1(\ram[103][5] ), .IN2(n458), .IN3(n549), .IN4(n222), .Q(
        n3249) );
  AO22X1 U1529 ( .IN1(\ram[103][6] ), .IN2(n458), .IN3(n549), .IN4(n255), .Q(
        n3250) );
  AO22X1 U1530 ( .IN1(\ram[103][7] ), .IN2(n458), .IN3(n549), .IN4(n288), .Q(
        n3251) );
  AO22X1 U1533 ( .IN1(\ram[102][0] ), .IN2(n461), .IN3(n4154), .IN4(n57), .Q(
        n3252) );
  AO22X1 U1534 ( .IN1(\ram[102][1] ), .IN2(n461), .IN3(n4154), .IN4(n90), .Q(
        n3253) );
  AO22X1 U1535 ( .IN1(\ram[102][2] ), .IN2(n461), .IN3(n4154), .IN4(n123), .Q(
        n3254) );
  AO22X1 U1536 ( .IN1(\ram[102][3] ), .IN2(n461), .IN3(n4154), .IN4(n156), .Q(
        n3255) );
  AO22X1 U1537 ( .IN1(\ram[102][4] ), .IN2(n461), .IN3(n4154), .IN4(n189), .Q(
        n3256) );
  AO22X1 U1538 ( .IN1(\ram[102][5] ), .IN2(n461), .IN3(n4154), .IN4(n222), .Q(
        n3257) );
  AO22X1 U1539 ( .IN1(\ram[102][6] ), .IN2(n461), .IN3(n4154), .IN4(n255), .Q(
        n3258) );
  AO22X1 U1540 ( .IN1(\ram[102][7] ), .IN2(n461), .IN3(n4154), .IN4(n288), .Q(
        n3259) );
  AO22X1 U1543 ( .IN1(\ram[101][0] ), .IN2(n464), .IN3(n645), .IN4(n57), .Q(
        n3260) );
  AO22X1 U1544 ( .IN1(\ram[101][1] ), .IN2(n464), .IN3(n645), .IN4(n90), .Q(
        n3261) );
  AO22X1 U1545 ( .IN1(\ram[101][2] ), .IN2(n464), .IN3(n645), .IN4(n123), .Q(
        n3262) );
  AO22X1 U1546 ( .IN1(\ram[101][3] ), .IN2(n464), .IN3(n645), .IN4(n156), .Q(
        n3263) );
  AO22X1 U1547 ( .IN1(\ram[101][4] ), .IN2(n464), .IN3(n645), .IN4(n189), .Q(
        n3264) );
  AO22X1 U1548 ( .IN1(\ram[101][5] ), .IN2(n464), .IN3(n645), .IN4(n222), .Q(
        n3265) );
  AO22X1 U1549 ( .IN1(\ram[101][6] ), .IN2(n464), .IN3(n645), .IN4(n255), .Q(
        n3266) );
  AO22X1 U1550 ( .IN1(\ram[101][7] ), .IN2(n464), .IN3(n645), .IN4(n288), .Q(
        n3267) );
  AO22X1 U1553 ( .IN1(\ram[100][0] ), .IN2(n467), .IN3(n4106), .IN4(n57), .Q(
        n3268) );
  AO22X1 U1554 ( .IN1(\ram[100][1] ), .IN2(n467), .IN3(n4106), .IN4(n90), .Q(
        n3269) );
  AO22X1 U1555 ( .IN1(\ram[100][2] ), .IN2(n467), .IN3(n4106), .IN4(n123), .Q(
        n3270) );
  AO22X1 U1556 ( .IN1(\ram[100][3] ), .IN2(n467), .IN3(n4106), .IN4(n156), .Q(
        n3271) );
  AO22X1 U1557 ( .IN1(\ram[100][4] ), .IN2(n467), .IN3(n4106), .IN4(n189), .Q(
        n3272) );
  AO22X1 U1558 ( .IN1(\ram[100][5] ), .IN2(n467), .IN3(n4106), .IN4(n222), .Q(
        n3273) );
  AO22X1 U1559 ( .IN1(\ram[100][6] ), .IN2(n467), .IN3(n4106), .IN4(n255), .Q(
        n3274) );
  AO22X1 U1560 ( .IN1(\ram[100][7] ), .IN2(n467), .IN3(n4106), .IN4(n288), .Q(
        n3275) );
  AO22X1 U1563 ( .IN1(\ram[99][0] ), .IN2(n470), .IN3(n501), .IN4(n57), .Q(
        n3276) );
  AO22X1 U1564 ( .IN1(\ram[99][1] ), .IN2(n470), .IN3(n501), .IN4(n90), .Q(
        n3277) );
  AO22X1 U1565 ( .IN1(\ram[99][2] ), .IN2(n470), .IN3(n501), .IN4(n123), .Q(
        n3278) );
  AO22X1 U1566 ( .IN1(\ram[99][3] ), .IN2(n470), .IN3(n501), .IN4(n156), .Q(
        n3279) );
  AO22X1 U1567 ( .IN1(\ram[99][4] ), .IN2(n470), .IN3(n501), .IN4(n189), .Q(
        n3280) );
  AO22X1 U1568 ( .IN1(\ram[99][5] ), .IN2(n470), .IN3(n501), .IN4(n222), .Q(
        n3281) );
  AO22X1 U1569 ( .IN1(\ram[99][6] ), .IN2(n470), .IN3(n501), .IN4(n255), .Q(
        n3282) );
  AO22X1 U1570 ( .IN1(\ram[99][7] ), .IN2(n470), .IN3(n501), .IN4(n288), .Q(
        n3283) );
  AO22X1 U1573 ( .IN1(\ram[98][0] ), .IN2(n473), .IN3(n4138), .IN4(n57), .Q(
        n3284) );
  AO22X1 U1574 ( .IN1(\ram[98][1] ), .IN2(n473), .IN3(n4138), .IN4(n90), .Q(
        n3285) );
  AO22X1 U1575 ( .IN1(\ram[98][2] ), .IN2(n473), .IN3(n4138), .IN4(n123), .Q(
        n3286) );
  AO22X1 U1576 ( .IN1(\ram[98][3] ), .IN2(n473), .IN3(n4138), .IN4(n156), .Q(
        n3287) );
  AO22X1 U1577 ( .IN1(\ram[98][4] ), .IN2(n473), .IN3(n4138), .IN4(n189), .Q(
        n3288) );
  AO22X1 U1578 ( .IN1(\ram[98][5] ), .IN2(n473), .IN3(n4138), .IN4(n222), .Q(
        n3289) );
  AO22X1 U1579 ( .IN1(\ram[98][6] ), .IN2(n473), .IN3(n4138), .IN4(n255), .Q(
        n3290) );
  AO22X1 U1580 ( .IN1(\ram[98][7] ), .IN2(n473), .IN3(n4138), .IN4(n288), .Q(
        n3291) );
  AO22X1 U1583 ( .IN1(\ram[97][0] ), .IN2(n476), .IN3(n597), .IN4(n57), .Q(
        n3292) );
  AO22X1 U1584 ( .IN1(\ram[97][1] ), .IN2(n476), .IN3(n597), .IN4(n90), .Q(
        n3293) );
  AO22X1 U1585 ( .IN1(\ram[97][2] ), .IN2(n476), .IN3(n597), .IN4(n123), .Q(
        n3294) );
  AO22X1 U1586 ( .IN1(\ram[97][3] ), .IN2(n476), .IN3(n597), .IN4(n156), .Q(
        n3295) );
  AO22X1 U1587 ( .IN1(\ram[97][4] ), .IN2(n476), .IN3(n597), .IN4(n189), .Q(
        n3296) );
  AO22X1 U1588 ( .IN1(\ram[97][5] ), .IN2(n476), .IN3(n597), .IN4(n222), .Q(
        n3297) );
  AO22X1 U1589 ( .IN1(\ram[97][6] ), .IN2(n476), .IN3(n597), .IN4(n255), .Q(
        n3298) );
  AO22X1 U1590 ( .IN1(\ram[97][7] ), .IN2(n476), .IN3(n597), .IN4(n288), .Q(
        n3299) );
  AO22X1 U1593 ( .IN1(\ram[96][0] ), .IN2(n479), .IN3(n4119), .IN4(n57), .Q(
        n3300) );
  AO22X1 U1594 ( .IN1(\ram[96][1] ), .IN2(n479), .IN3(n4119), .IN4(n90), .Q(
        n3301) );
  AO22X1 U1595 ( .IN1(\ram[96][2] ), .IN2(n479), .IN3(n4119), .IN4(n123), .Q(
        n3302) );
  AO22X1 U1596 ( .IN1(\ram[96][3] ), .IN2(n479), .IN3(n4119), .IN4(n156), .Q(
        n3303) );
  AO22X1 U1597 ( .IN1(\ram[96][4] ), .IN2(n479), .IN3(n4119), .IN4(n189), .Q(
        n3304) );
  AO22X1 U1598 ( .IN1(\ram[96][5] ), .IN2(n479), .IN3(n4119), .IN4(n222), .Q(
        n3305) );
  AO22X1 U1599 ( .IN1(\ram[96][6] ), .IN2(n479), .IN3(n4119), .IN4(n255), .Q(
        n3306) );
  AO22X1 U1600 ( .IN1(\ram[96][7] ), .IN2(n479), .IN3(n4119), .IN4(n288), .Q(
        n3307) );
  AO22X1 U1603 ( .IN1(\ram[95][0] ), .IN2(n482), .IN3(n348), .IN4(n54), .Q(
        n3308) );
  AO22X1 U1604 ( .IN1(\ram[95][1] ), .IN2(n482), .IN3(n348), .IN4(n87), .Q(
        n3309) );
  AO22X1 U1605 ( .IN1(\ram[95][2] ), .IN2(n482), .IN3(n348), .IN4(n120), .Q(
        n3310) );
  AO22X1 U1606 ( .IN1(\ram[95][3] ), .IN2(n482), .IN3(n348), .IN4(n153), .Q(
        n3311) );
  AO22X1 U1607 ( .IN1(\ram[95][4] ), .IN2(n482), .IN3(n348), .IN4(n186), .Q(
        n3312) );
  AO22X1 U1608 ( .IN1(\ram[95][5] ), .IN2(n482), .IN3(n348), .IN4(n219), .Q(
        n3313) );
  AO22X1 U1609 ( .IN1(\ram[95][6] ), .IN2(n482), .IN3(n348), .IN4(n252), .Q(
        n3314) );
  AO22X1 U1610 ( .IN1(\ram[95][7] ), .IN2(n482), .IN3(n348), .IN4(n285), .Q(
        n3315) );
  AO22X1 U1613 ( .IN1(\ram[94][0] ), .IN2(n485), .IN3(n4090), .IN4(n54), .Q(
        n3316) );
  AO22X1 U1614 ( .IN1(\ram[94][1] ), .IN2(n485), .IN3(n4090), .IN4(n87), .Q(
        n3317) );
  AO22X1 U1615 ( .IN1(\ram[94][2] ), .IN2(n485), .IN3(n4090), .IN4(n120), .Q(
        n3318) );
  AO22X1 U1616 ( .IN1(\ram[94][3] ), .IN2(n485), .IN3(n4090), .IN4(n153), .Q(
        n3319) );
  AO22X1 U1617 ( .IN1(\ram[94][4] ), .IN2(n485), .IN3(n4090), .IN4(n186), .Q(
        n3320) );
  AO22X1 U1618 ( .IN1(\ram[94][5] ), .IN2(n485), .IN3(n4090), .IN4(n219), .Q(
        n3321) );
  AO22X1 U1619 ( .IN1(\ram[94][6] ), .IN2(n485), .IN3(n4090), .IN4(n252), .Q(
        n3322) );
  AO22X1 U1620 ( .IN1(\ram[94][7] ), .IN2(n485), .IN3(n4090), .IN4(n285), .Q(
        n3323) );
  AO22X1 U1623 ( .IN1(\ram[93][0] ), .IN2(n488), .IN3(n453), .IN4(n54), .Q(
        n3324) );
  AO22X1 U1624 ( .IN1(\ram[93][1] ), .IN2(n488), .IN3(n453), .IN4(n87), .Q(
        n3325) );
  AO22X1 U1625 ( .IN1(\ram[93][2] ), .IN2(n488), .IN3(n453), .IN4(n120), .Q(
        n3326) );
  AO22X1 U1626 ( .IN1(\ram[93][3] ), .IN2(n488), .IN3(n453), .IN4(n153), .Q(
        n3327) );
  AO22X1 U1627 ( .IN1(\ram[93][4] ), .IN2(n488), .IN3(n453), .IN4(n186), .Q(
        n3328) );
  AO22X1 U1628 ( .IN1(\ram[93][5] ), .IN2(n488), .IN3(n453), .IN4(n219), .Q(
        n3329) );
  AO22X1 U1629 ( .IN1(\ram[93][6] ), .IN2(n488), .IN3(n453), .IN4(n252), .Q(
        n3330) );
  AO22X1 U1630 ( .IN1(\ram[93][7] ), .IN2(n488), .IN3(n453), .IN4(n285), .Q(
        n3331) );
  AO22X1 U1633 ( .IN1(\ram[92][0] ), .IN2(n491), .IN3(n735), .IN4(n54), .Q(
        n3332) );
  AO22X1 U1634 ( .IN1(\ram[92][1] ), .IN2(n491), .IN3(n735), .IN4(n87), .Q(
        n3333) );
  AO22X1 U1635 ( .IN1(\ram[92][2] ), .IN2(n491), .IN3(n735), .IN4(n120), .Q(
        n3334) );
  AO22X1 U1636 ( .IN1(\ram[92][3] ), .IN2(n491), .IN3(n735), .IN4(n153), .Q(
        n3335) );
  AO22X1 U1637 ( .IN1(\ram[92][4] ), .IN2(n491), .IN3(n735), .IN4(n186), .Q(
        n3336) );
  AO22X1 U1638 ( .IN1(\ram[92][5] ), .IN2(n491), .IN3(n735), .IN4(n219), .Q(
        n3337) );
  AO22X1 U1639 ( .IN1(\ram[92][6] ), .IN2(n491), .IN3(n735), .IN4(n252), .Q(
        n3338) );
  AO22X1 U1640 ( .IN1(\ram[92][7] ), .IN2(n491), .IN3(n735), .IN4(n285), .Q(
        n3339) );
  AO22X1 U1643 ( .IN1(\ram[91][0] ), .IN2(n494), .IN3(n300), .IN4(n54), .Q(
        n3340) );
  AO22X1 U1644 ( .IN1(\ram[91][1] ), .IN2(n494), .IN3(n300), .IN4(n87), .Q(
        n3341) );
  AO22X1 U1645 ( .IN1(\ram[91][2] ), .IN2(n494), .IN3(n300), .IN4(n120), .Q(
        n3342) );
  AO22X1 U1646 ( .IN1(\ram[91][3] ), .IN2(n494), .IN3(n300), .IN4(n153), .Q(
        n3343) );
  AO22X1 U1647 ( .IN1(\ram[91][4] ), .IN2(n494), .IN3(n300), .IN4(n186), .Q(
        n3344) );
  AO22X1 U1648 ( .IN1(\ram[91][5] ), .IN2(n494), .IN3(n300), .IN4(n219), .Q(
        n3345) );
  AO22X1 U1649 ( .IN1(\ram[91][6] ), .IN2(n494), .IN3(n300), .IN4(n252), .Q(
        n3346) );
  AO22X1 U1650 ( .IN1(\ram[91][7] ), .IN2(n494), .IN3(n300), .IN4(n285), .Q(
        n3347) );
  AO22X1 U1653 ( .IN1(\ram[90][0] ), .IN2(n497), .IN3(n2015), .IN4(n54), .Q(
        n3348) );
  AO22X1 U1654 ( .IN1(\ram[90][1] ), .IN2(n497), .IN3(n2015), .IN4(n87), .Q(
        n3349) );
  AO22X1 U1655 ( .IN1(\ram[90][2] ), .IN2(n497), .IN3(n2015), .IN4(n120), .Q(
        n3350) );
  AO22X1 U1656 ( .IN1(\ram[90][3] ), .IN2(n497), .IN3(n2015), .IN4(n153), .Q(
        n3351) );
  AO22X1 U1657 ( .IN1(\ram[90][4] ), .IN2(n497), .IN3(n2015), .IN4(n186), .Q(
        n3352) );
  AO22X1 U1658 ( .IN1(\ram[90][5] ), .IN2(n497), .IN3(n2015), .IN4(n219), .Q(
        n3353) );
  AO22X1 U1659 ( .IN1(\ram[90][6] ), .IN2(n497), .IN3(n2015), .IN4(n252), .Q(
        n3354) );
  AO22X1 U1660 ( .IN1(\ram[90][7] ), .IN2(n497), .IN3(n2015), .IN4(n285), .Q(
        n3355) );
  AO22X1 U1663 ( .IN1(\ram[89][0] ), .IN2(n500), .IN3(n399), .IN4(n54), .Q(
        n3356) );
  AO22X1 U1664 ( .IN1(\ram[89][1] ), .IN2(n500), .IN3(n399), .IN4(n87), .Q(
        n3357) );
  AO22X1 U1665 ( .IN1(\ram[89][2] ), .IN2(n500), .IN3(n399), .IN4(n120), .Q(
        n3358) );
  AO22X1 U1666 ( .IN1(\ram[89][3] ), .IN2(n500), .IN3(n399), .IN4(n153), .Q(
        n3359) );
  AO22X1 U1667 ( .IN1(\ram[89][4] ), .IN2(n500), .IN3(n399), .IN4(n186), .Q(
        n3360) );
  AO22X1 U1668 ( .IN1(\ram[89][5] ), .IN2(n500), .IN3(n399), .IN4(n219), .Q(
        n3361) );
  AO22X1 U1669 ( .IN1(\ram[89][6] ), .IN2(n500), .IN3(n399), .IN4(n252), .Q(
        n3362) );
  AO22X1 U1670 ( .IN1(\ram[89][7] ), .IN2(n500), .IN3(n399), .IN4(n285), .Q(
        n3363) );
  AO22X1 U1673 ( .IN1(\ram[88][0] ), .IN2(n503), .IN3(n687), .IN4(n54), .Q(
        n3364) );
  AO22X1 U1674 ( .IN1(\ram[88][1] ), .IN2(n503), .IN3(n687), .IN4(n87), .Q(
        n3365) );
  AO22X1 U1675 ( .IN1(\ram[88][2] ), .IN2(n503), .IN3(n687), .IN4(n120), .Q(
        n3366) );
  AO22X1 U1676 ( .IN1(\ram[88][3] ), .IN2(n503), .IN3(n687), .IN4(n153), .Q(
        n3367) );
  AO22X1 U1677 ( .IN1(\ram[88][4] ), .IN2(n503), .IN3(n687), .IN4(n186), .Q(
        n3368) );
  AO22X1 U1678 ( .IN1(\ram[88][5] ), .IN2(n503), .IN3(n687), .IN4(n219), .Q(
        n3369) );
  AO22X1 U1679 ( .IN1(\ram[88][6] ), .IN2(n503), .IN3(n687), .IN4(n252), .Q(
        n3370) );
  AO22X1 U1680 ( .IN1(\ram[88][7] ), .IN2(n503), .IN3(n687), .IN4(n285), .Q(
        n3371) );
  AO22X1 U1683 ( .IN1(\ram[87][0] ), .IN2(n506), .IN3(n540), .IN4(n54), .Q(
        n3372) );
  AO22X1 U1684 ( .IN1(\ram[87][1] ), .IN2(n506), .IN3(n540), .IN4(n87), .Q(
        n3373) );
  AO22X1 U1685 ( .IN1(\ram[87][2] ), .IN2(n506), .IN3(n540), .IN4(n120), .Q(
        n3374) );
  AO22X1 U1686 ( .IN1(\ram[87][3] ), .IN2(n506), .IN3(n540), .IN4(n153), .Q(
        n3375) );
  AO22X1 U1687 ( .IN1(\ram[87][4] ), .IN2(n506), .IN3(n540), .IN4(n186), .Q(
        n3376) );
  AO22X1 U1688 ( .IN1(\ram[87][5] ), .IN2(n506), .IN3(n540), .IN4(n219), .Q(
        n3377) );
  AO22X1 U1689 ( .IN1(\ram[87][6] ), .IN2(n506), .IN3(n540), .IN4(n252), .Q(
        n3378) );
  AO22X1 U1690 ( .IN1(\ram[87][7] ), .IN2(n506), .IN3(n540), .IN4(n285), .Q(
        n3379) );
  AO22X1 U1693 ( .IN1(\ram[86][0] ), .IN2(n509), .IN3(n4151), .IN4(n54), .Q(
        n3380) );
  AO22X1 U1694 ( .IN1(\ram[86][1] ), .IN2(n509), .IN3(n4151), .IN4(n87), .Q(
        n3381) );
  AO22X1 U1695 ( .IN1(\ram[86][2] ), .IN2(n509), .IN3(n4151), .IN4(n120), .Q(
        n3382) );
  AO22X1 U1696 ( .IN1(\ram[86][3] ), .IN2(n509), .IN3(n4151), .IN4(n153), .Q(
        n3383) );
  AO22X1 U1697 ( .IN1(\ram[86][4] ), .IN2(n509), .IN3(n4151), .IN4(n186), .Q(
        n3384) );
  AO22X1 U1698 ( .IN1(\ram[86][5] ), .IN2(n509), .IN3(n4151), .IN4(n219), .Q(
        n3385) );
  AO22X1 U1699 ( .IN1(\ram[86][6] ), .IN2(n509), .IN3(n4151), .IN4(n252), .Q(
        n3386) );
  AO22X1 U1700 ( .IN1(\ram[86][7] ), .IN2(n509), .IN3(n4151), .IN4(n285), .Q(
        n3387) );
  AO22X1 U1703 ( .IN1(\ram[85][0] ), .IN2(n512), .IN3(n636), .IN4(n54), .Q(
        n3388) );
  AO22X1 U1704 ( .IN1(\ram[85][1] ), .IN2(n512), .IN3(n636), .IN4(n87), .Q(
        n3389) );
  AO22X1 U1705 ( .IN1(\ram[85][2] ), .IN2(n512), .IN3(n636), .IN4(n120), .Q(
        n3390) );
  AO22X1 U1706 ( .IN1(\ram[85][3] ), .IN2(n512), .IN3(n636), .IN4(n153), .Q(
        n3391) );
  AO22X1 U1707 ( .IN1(\ram[85][4] ), .IN2(n512), .IN3(n636), .IN4(n186), .Q(
        n3392) );
  AO22X1 U1708 ( .IN1(\ram[85][5] ), .IN2(n512), .IN3(n636), .IN4(n219), .Q(
        n3393) );
  AO22X1 U1709 ( .IN1(\ram[85][6] ), .IN2(n512), .IN3(n636), .IN4(n252), .Q(
        n3394) );
  AO22X1 U1710 ( .IN1(\ram[85][7] ), .IN2(n512), .IN3(n636), .IN4(n285), .Q(
        n3395) );
  AO22X1 U1713 ( .IN1(\ram[84][0] ), .IN2(n515), .IN3(n4103), .IN4(n54), .Q(
        n3396) );
  AO22X1 U1714 ( .IN1(\ram[84][1] ), .IN2(n515), .IN3(n4103), .IN4(n87), .Q(
        n3397) );
  AO22X1 U1715 ( .IN1(\ram[84][2] ), .IN2(n515), .IN3(n4103), .IN4(n120), .Q(
        n3398) );
  AO22X1 U1716 ( .IN1(\ram[84][3] ), .IN2(n515), .IN3(n4103), .IN4(n153), .Q(
        n3399) );
  AO22X1 U1717 ( .IN1(\ram[84][4] ), .IN2(n515), .IN3(n4103), .IN4(n186), .Q(
        n3400) );
  AO22X1 U1718 ( .IN1(\ram[84][5] ), .IN2(n515), .IN3(n4103), .IN4(n219), .Q(
        n3401) );
  AO22X1 U1719 ( .IN1(\ram[84][6] ), .IN2(n515), .IN3(n4103), .IN4(n252), .Q(
        n3402) );
  AO22X1 U1720 ( .IN1(\ram[84][7] ), .IN2(n515), .IN3(n4103), .IN4(n285), .Q(
        n3403) );
  AO22X1 U1723 ( .IN1(\ram[83][0] ), .IN2(n518), .IN3(n492), .IN4(datain[0]), 
        .Q(n3404) );
  AO22X1 U1724 ( .IN1(\ram[83][1] ), .IN2(n518), .IN3(n492), .IN4(datain[1]), 
        .Q(n3405) );
  AO22X1 U1725 ( .IN1(\ram[83][2] ), .IN2(n518), .IN3(n492), .IN4(datain[2]), 
        .Q(n3406) );
  AO22X1 U1726 ( .IN1(\ram[83][3] ), .IN2(n518), .IN3(n492), .IN4(datain[3]), 
        .Q(n3407) );
  AO22X1 U1727 ( .IN1(\ram[83][4] ), .IN2(n518), .IN3(n492), .IN4(datain[4]), 
        .Q(n3408) );
  AO22X1 U1728 ( .IN1(\ram[83][5] ), .IN2(n518), .IN3(n492), .IN4(datain[5]), 
        .Q(n3409) );
  AO22X1 U1729 ( .IN1(\ram[83][6] ), .IN2(n518), .IN3(n492), .IN4(datain[6]), 
        .Q(n3410) );
  AO22X1 U1730 ( .IN1(\ram[83][7] ), .IN2(n518), .IN3(n492), .IN4(datain[7]), 
        .Q(n3411) );
  AO22X1 U1733 ( .IN1(\ram[82][0] ), .IN2(n521), .IN3(n4135), .IN4(datain[0]), 
        .Q(n3412) );
  AO22X1 U1734 ( .IN1(\ram[82][1] ), .IN2(n521), .IN3(n4135), .IN4(datain[1]), 
        .Q(n3413) );
  AO22X1 U1735 ( .IN1(\ram[82][2] ), .IN2(n521), .IN3(n4135), .IN4(datain[2]), 
        .Q(n3414) );
  AO22X1 U1736 ( .IN1(\ram[82][3] ), .IN2(n521), .IN3(n4135), .IN4(datain[3]), 
        .Q(n3415) );
  AO22X1 U1737 ( .IN1(\ram[82][4] ), .IN2(n521), .IN3(n4135), .IN4(datain[4]), 
        .Q(n3416) );
  AO22X1 U1738 ( .IN1(\ram[82][5] ), .IN2(n521), .IN3(n4135), .IN4(datain[5]), 
        .Q(n3417) );
  AO22X1 U1739 ( .IN1(\ram[82][6] ), .IN2(n521), .IN3(n4135), .IN4(datain[6]), 
        .Q(n3418) );
  AO22X1 U1740 ( .IN1(\ram[82][7] ), .IN2(n521), .IN3(n4135), .IN4(datain[7]), 
        .Q(n3419) );
  AO22X1 U1743 ( .IN1(\ram[81][0] ), .IN2(n524), .IN3(n588), .IN4(datain[0]), 
        .Q(n3420) );
  AO22X1 U1744 ( .IN1(\ram[81][1] ), .IN2(n524), .IN3(n588), .IN4(datain[1]), 
        .Q(n3421) );
  AO22X1 U1745 ( .IN1(\ram[81][2] ), .IN2(n524), .IN3(n588), .IN4(datain[2]), 
        .Q(n3422) );
  AO22X1 U1746 ( .IN1(\ram[81][3] ), .IN2(n524), .IN3(n588), .IN4(datain[3]), 
        .Q(n3423) );
  AO22X1 U1747 ( .IN1(\ram[81][4] ), .IN2(n524), .IN3(n588), .IN4(datain[4]), 
        .Q(n3424) );
  AO22X1 U1748 ( .IN1(\ram[81][5] ), .IN2(n524), .IN3(n588), .IN4(datain[5]), 
        .Q(n3425) );
  AO22X1 U1749 ( .IN1(\ram[81][6] ), .IN2(n524), .IN3(n588), .IN4(datain[6]), 
        .Q(n3426) );
  AO22X1 U1750 ( .IN1(\ram[81][7] ), .IN2(n524), .IN3(n588), .IN4(datain[7]), 
        .Q(n3427) );
  AO22X1 U1753 ( .IN1(\ram[80][0] ), .IN2(n527), .IN3(n4120), .IN4(datain[0]), 
        .Q(n3428) );
  AO22X1 U1754 ( .IN1(\ram[80][1] ), .IN2(n527), .IN3(n4120), .IN4(datain[1]), 
        .Q(n3429) );
  AO22X1 U1755 ( .IN1(\ram[80][2] ), .IN2(n527), .IN3(n4120), .IN4(datain[2]), 
        .Q(n3430) );
  AO22X1 U1756 ( .IN1(\ram[80][3] ), .IN2(n527), .IN3(n4120), .IN4(datain[3]), 
        .Q(n3431) );
  AO22X1 U1757 ( .IN1(\ram[80][4] ), .IN2(n527), .IN3(n4120), .IN4(datain[4]), 
        .Q(n3432) );
  AO22X1 U1758 ( .IN1(\ram[80][5] ), .IN2(n527), .IN3(n4120), .IN4(datain[5]), 
        .Q(n3433) );
  AO22X1 U1759 ( .IN1(\ram[80][6] ), .IN2(n527), .IN3(n4120), .IN4(datain[6]), 
        .Q(n3434) );
  AO22X1 U1760 ( .IN1(\ram[80][7] ), .IN2(n527), .IN3(n4120), .IN4(datain[7]), 
        .Q(n3435) );
  AO22X1 U1763 ( .IN1(\ram[79][0] ), .IN2(n530), .IN3(n351), .IN4(datain[0]), 
        .Q(n3436) );
  AO22X1 U1764 ( .IN1(\ram[79][1] ), .IN2(n530), .IN3(n351), .IN4(datain[1]), 
        .Q(n3437) );
  AO22X1 U1765 ( .IN1(\ram[79][2] ), .IN2(n530), .IN3(n351), .IN4(datain[2]), 
        .Q(n3438) );
  AO22X1 U1766 ( .IN1(\ram[79][3] ), .IN2(n530), .IN3(n351), .IN4(datain[3]), 
        .Q(n3439) );
  AO22X1 U1767 ( .IN1(\ram[79][4] ), .IN2(n530), .IN3(n351), .IN4(datain[4]), 
        .Q(n3440) );
  AO22X1 U1768 ( .IN1(\ram[79][5] ), .IN2(n530), .IN3(n351), .IN4(datain[5]), 
        .Q(n3441) );
  AO22X1 U1769 ( .IN1(\ram[79][6] ), .IN2(n530), .IN3(n351), .IN4(datain[6]), 
        .Q(n3442) );
  AO22X1 U1770 ( .IN1(\ram[79][7] ), .IN2(n530), .IN3(n351), .IN4(datain[7]), 
        .Q(n3443) );
  AO22X1 U1773 ( .IN1(\ram[78][0] ), .IN2(n533), .IN3(n4091), .IN4(datain[0]), 
        .Q(n3444) );
  AO22X1 U1774 ( .IN1(\ram[78][1] ), .IN2(n533), .IN3(n4091), .IN4(datain[1]), 
        .Q(n3445) );
  AO22X1 U1775 ( .IN1(\ram[78][2] ), .IN2(n533), .IN3(n4091), .IN4(datain[2]), 
        .Q(n3446) );
  AO22X1 U1776 ( .IN1(\ram[78][3] ), .IN2(n533), .IN3(n4091), .IN4(datain[3]), 
        .Q(n3447) );
  AO22X1 U1777 ( .IN1(\ram[78][4] ), .IN2(n533), .IN3(n4091), .IN4(datain[4]), 
        .Q(n3448) );
  AO22X1 U1778 ( .IN1(\ram[78][5] ), .IN2(n533), .IN3(n4091), .IN4(datain[5]), 
        .Q(n3449) );
  AO22X1 U1779 ( .IN1(\ram[78][6] ), .IN2(n533), .IN3(n4091), .IN4(datain[6]), 
        .Q(n3450) );
  AO22X1 U1780 ( .IN1(\ram[78][7] ), .IN2(n533), .IN3(n4091), .IN4(datain[7]), 
        .Q(n3451) );
  AO22X1 U1783 ( .IN1(\ram[77][0] ), .IN2(n536), .IN3(n456), .IN4(datain[0]), 
        .Q(n3452) );
  AO22X1 U1784 ( .IN1(\ram[77][1] ), .IN2(n536), .IN3(n456), .IN4(datain[1]), 
        .Q(n3453) );
  AO22X1 U1785 ( .IN1(\ram[77][2] ), .IN2(n536), .IN3(n456), .IN4(datain[2]), 
        .Q(n3454) );
  AO22X1 U1786 ( .IN1(\ram[77][3] ), .IN2(n536), .IN3(n456), .IN4(datain[3]), 
        .Q(n3455) );
  AO22X1 U1787 ( .IN1(\ram[77][4] ), .IN2(n536), .IN3(n456), .IN4(datain[4]), 
        .Q(n3456) );
  AO22X1 U1788 ( .IN1(\ram[77][5] ), .IN2(n536), .IN3(n456), .IN4(datain[5]), 
        .Q(n3457) );
  AO22X1 U1789 ( .IN1(\ram[77][6] ), .IN2(n536), .IN3(n456), .IN4(datain[6]), 
        .Q(n3458) );
  AO22X1 U1790 ( .IN1(\ram[77][7] ), .IN2(n536), .IN3(n456), .IN4(datain[7]), 
        .Q(n3459) );
  AO22X1 U1793 ( .IN1(\ram[76][0] ), .IN2(n539), .IN3(n738), .IN4(datain[0]), 
        .Q(n3460) );
  AO22X1 U1794 ( .IN1(\ram[76][1] ), .IN2(n539), .IN3(n738), .IN4(datain[1]), 
        .Q(n3461) );
  AO22X1 U1795 ( .IN1(\ram[76][2] ), .IN2(n539), .IN3(n738), .IN4(datain[2]), 
        .Q(n3462) );
  AO22X1 U1796 ( .IN1(\ram[76][3] ), .IN2(n539), .IN3(n738), .IN4(datain[3]), 
        .Q(n3463) );
  AO22X1 U1797 ( .IN1(\ram[76][4] ), .IN2(n539), .IN3(n738), .IN4(datain[4]), 
        .Q(n3464) );
  AO22X1 U1798 ( .IN1(\ram[76][5] ), .IN2(n539), .IN3(n738), .IN4(datain[5]), 
        .Q(n3465) );
  AO22X1 U1799 ( .IN1(\ram[76][6] ), .IN2(n539), .IN3(n738), .IN4(datain[6]), 
        .Q(n3466) );
  AO22X1 U1800 ( .IN1(\ram[76][7] ), .IN2(n539), .IN3(n738), .IN4(datain[7]), 
        .Q(n3467) );
  AO22X1 U1803 ( .IN1(\ram[75][0] ), .IN2(n542), .IN3(n303), .IN4(datain[0]), 
        .Q(n3468) );
  AO22X1 U1804 ( .IN1(\ram[75][1] ), .IN2(n542), .IN3(n303), .IN4(datain[1]), 
        .Q(n3469) );
  AO22X1 U1805 ( .IN1(\ram[75][2] ), .IN2(n542), .IN3(n303), .IN4(datain[2]), 
        .Q(n3470) );
  AO22X1 U1806 ( .IN1(\ram[75][3] ), .IN2(n542), .IN3(n303), .IN4(datain[3]), 
        .Q(n3471) );
  AO22X1 U1807 ( .IN1(\ram[75][4] ), .IN2(n542), .IN3(n303), .IN4(datain[4]), 
        .Q(n3472) );
  AO22X1 U1808 ( .IN1(\ram[75][5] ), .IN2(n542), .IN3(n303), .IN4(datain[5]), 
        .Q(n3473) );
  AO22X1 U1809 ( .IN1(\ram[75][6] ), .IN2(n542), .IN3(n303), .IN4(datain[6]), 
        .Q(n3474) );
  AO22X1 U1810 ( .IN1(\ram[75][7] ), .IN2(n542), .IN3(n303), .IN4(datain[7]), 
        .Q(n3475) );
  AO22X1 U1813 ( .IN1(\ram[74][0] ), .IN2(n545), .IN3(n2016), .IN4(datain[0]), 
        .Q(n3476) );
  AO22X1 U1814 ( .IN1(\ram[74][1] ), .IN2(n545), .IN3(n2016), .IN4(datain[1]), 
        .Q(n3477) );
  AO22X1 U1815 ( .IN1(\ram[74][2] ), .IN2(n545), .IN3(n2016), .IN4(datain[2]), 
        .Q(n3478) );
  AO22X1 U1816 ( .IN1(\ram[74][3] ), .IN2(n545), .IN3(n2016), .IN4(datain[3]), 
        .Q(n3479) );
  AO22X1 U1817 ( .IN1(\ram[74][4] ), .IN2(n545), .IN3(n2016), .IN4(datain[4]), 
        .Q(n3480) );
  AO22X1 U1818 ( .IN1(\ram[74][5] ), .IN2(n545), .IN3(n2016), .IN4(datain[5]), 
        .Q(n3481) );
  AO22X1 U1819 ( .IN1(\ram[74][6] ), .IN2(n545), .IN3(n2016), .IN4(datain[6]), 
        .Q(n3482) );
  AO22X1 U1820 ( .IN1(\ram[74][7] ), .IN2(n545), .IN3(n2016), .IN4(datain[7]), 
        .Q(n3483) );
  AO22X1 U1823 ( .IN1(\ram[73][0] ), .IN2(n548), .IN3(n402), .IN4(datain[0]), 
        .Q(n3484) );
  AO22X1 U1824 ( .IN1(\ram[73][1] ), .IN2(n548), .IN3(n402), .IN4(datain[1]), 
        .Q(n3485) );
  AO22X1 U1825 ( .IN1(\ram[73][2] ), .IN2(n548), .IN3(n402), .IN4(datain[2]), 
        .Q(n3486) );
  AO22X1 U1826 ( .IN1(\ram[73][3] ), .IN2(n548), .IN3(n402), .IN4(datain[3]), 
        .Q(n3487) );
  AO22X1 U1827 ( .IN1(\ram[73][4] ), .IN2(n548), .IN3(n402), .IN4(datain[4]), 
        .Q(n3488) );
  AO22X1 U1828 ( .IN1(\ram[73][5] ), .IN2(n548), .IN3(n402), .IN4(datain[5]), 
        .Q(n3489) );
  AO22X1 U1829 ( .IN1(\ram[73][6] ), .IN2(n548), .IN3(n402), .IN4(datain[6]), 
        .Q(n3490) );
  AO22X1 U1830 ( .IN1(\ram[73][7] ), .IN2(n548), .IN3(n402), .IN4(datain[7]), 
        .Q(n3491) );
  AO22X1 U1833 ( .IN1(\ram[72][0] ), .IN2(n551), .IN3(n690), .IN4(datain[0]), 
        .Q(n3492) );
  AO22X1 U1834 ( .IN1(\ram[72][1] ), .IN2(n551), .IN3(n690), .IN4(datain[1]), 
        .Q(n3493) );
  AO22X1 U1835 ( .IN1(\ram[72][2] ), .IN2(n551), .IN3(n690), .IN4(datain[2]), 
        .Q(n3494) );
  AO22X1 U1836 ( .IN1(\ram[72][3] ), .IN2(n551), .IN3(n690), .IN4(datain[3]), 
        .Q(n3495) );
  AO22X1 U1837 ( .IN1(\ram[72][4] ), .IN2(n551), .IN3(n690), .IN4(datain[4]), 
        .Q(n3496) );
  AO22X1 U1838 ( .IN1(\ram[72][5] ), .IN2(n551), .IN3(n690), .IN4(datain[5]), 
        .Q(n3497) );
  AO22X1 U1839 ( .IN1(\ram[72][6] ), .IN2(n551), .IN3(n690), .IN4(datain[6]), 
        .Q(n3498) );
  AO22X1 U1840 ( .IN1(\ram[72][7] ), .IN2(n551), .IN3(n690), .IN4(datain[7]), 
        .Q(n3499) );
  AO22X1 U1843 ( .IN1(\ram[71][0] ), .IN2(n554), .IN3(n543), .IN4(n51), .Q(
        n3500) );
  AO22X1 U1844 ( .IN1(\ram[71][1] ), .IN2(n554), .IN3(n543), .IN4(n84), .Q(
        n3501) );
  AO22X1 U1845 ( .IN1(\ram[71][2] ), .IN2(n554), .IN3(n543), .IN4(n117), .Q(
        n3502) );
  AO22X1 U1846 ( .IN1(\ram[71][3] ), .IN2(n554), .IN3(n543), .IN4(n150), .Q(
        n3503) );
  AO22X1 U1847 ( .IN1(\ram[71][4] ), .IN2(n554), .IN3(n543), .IN4(n183), .Q(
        n3504) );
  AO22X1 U1848 ( .IN1(\ram[71][5] ), .IN2(n554), .IN3(n543), .IN4(n216), .Q(
        n3505) );
  AO22X1 U1849 ( .IN1(\ram[71][6] ), .IN2(n554), .IN3(n543), .IN4(n249), .Q(
        n3506) );
  AO22X1 U1850 ( .IN1(\ram[71][7] ), .IN2(n554), .IN3(n543), .IN4(n282), .Q(
        n3507) );
  AO22X1 U1853 ( .IN1(\ram[70][0] ), .IN2(n557), .IN3(n4152), .IN4(n51), .Q(
        n3508) );
  AO22X1 U1854 ( .IN1(\ram[70][1] ), .IN2(n557), .IN3(n4152), .IN4(n84), .Q(
        n3509) );
  AO22X1 U1855 ( .IN1(\ram[70][2] ), .IN2(n557), .IN3(n4152), .IN4(n117), .Q(
        n3510) );
  AO22X1 U1856 ( .IN1(\ram[70][3] ), .IN2(n557), .IN3(n4152), .IN4(n150), .Q(
        n3511) );
  AO22X1 U1857 ( .IN1(\ram[70][4] ), .IN2(n557), .IN3(n4152), .IN4(n183), .Q(
        n3512) );
  AO22X1 U1858 ( .IN1(\ram[70][5] ), .IN2(n557), .IN3(n4152), .IN4(n216), .Q(
        n3513) );
  AO22X1 U1859 ( .IN1(\ram[70][6] ), .IN2(n557), .IN3(n4152), .IN4(n249), .Q(
        n3514) );
  AO22X1 U1860 ( .IN1(\ram[70][7] ), .IN2(n557), .IN3(n4152), .IN4(n282), .Q(
        n3515) );
  AO22X1 U1863 ( .IN1(\ram[69][0] ), .IN2(n560), .IN3(n639), .IN4(n51), .Q(
        n3516) );
  AO22X1 U1864 ( .IN1(\ram[69][1] ), .IN2(n560), .IN3(n639), .IN4(n84), .Q(
        n3517) );
  AO22X1 U1865 ( .IN1(\ram[69][2] ), .IN2(n560), .IN3(n639), .IN4(n117), .Q(
        n3518) );
  AO22X1 U1866 ( .IN1(\ram[69][3] ), .IN2(n560), .IN3(n639), .IN4(n150), .Q(
        n3519) );
  AO22X1 U1867 ( .IN1(\ram[69][4] ), .IN2(n560), .IN3(n639), .IN4(n183), .Q(
        n3520) );
  AO22X1 U1868 ( .IN1(\ram[69][5] ), .IN2(n560), .IN3(n639), .IN4(n216), .Q(
        n3521) );
  AO22X1 U1869 ( .IN1(\ram[69][6] ), .IN2(n560), .IN3(n639), .IN4(n249), .Q(
        n3522) );
  AO22X1 U1870 ( .IN1(\ram[69][7] ), .IN2(n560), .IN3(n639), .IN4(n282), .Q(
        n3523) );
  AO22X1 U1873 ( .IN1(\ram[68][0] ), .IN2(n563), .IN3(n4104), .IN4(n51), .Q(
        n3524) );
  AO22X1 U1874 ( .IN1(\ram[68][1] ), .IN2(n563), .IN3(n4104), .IN4(n84), .Q(
        n3525) );
  AO22X1 U1875 ( .IN1(\ram[68][2] ), .IN2(n563), .IN3(n4104), .IN4(n117), .Q(
        n3526) );
  AO22X1 U1876 ( .IN1(\ram[68][3] ), .IN2(n563), .IN3(n4104), .IN4(n150), .Q(
        n3527) );
  AO22X1 U1877 ( .IN1(\ram[68][4] ), .IN2(n563), .IN3(n4104), .IN4(n183), .Q(
        n3528) );
  AO22X1 U1878 ( .IN1(\ram[68][5] ), .IN2(n563), .IN3(n4104), .IN4(n216), .Q(
        n3529) );
  AO22X1 U1879 ( .IN1(\ram[68][6] ), .IN2(n563), .IN3(n4104), .IN4(n249), .Q(
        n3530) );
  AO22X1 U1880 ( .IN1(\ram[68][7] ), .IN2(n563), .IN3(n4104), .IN4(n282), .Q(
        n3531) );
  AO22X1 U1883 ( .IN1(\ram[67][0] ), .IN2(n566), .IN3(n495), .IN4(n51), .Q(
        n3532) );
  AO22X1 U1884 ( .IN1(\ram[67][1] ), .IN2(n566), .IN3(n495), .IN4(n84), .Q(
        n3533) );
  AO22X1 U1885 ( .IN1(\ram[67][2] ), .IN2(n566), .IN3(n495), .IN4(n117), .Q(
        n3534) );
  AO22X1 U1886 ( .IN1(\ram[67][3] ), .IN2(n566), .IN3(n495), .IN4(n150), .Q(
        n3535) );
  AO22X1 U1887 ( .IN1(\ram[67][4] ), .IN2(n566), .IN3(n495), .IN4(n183), .Q(
        n3536) );
  AO22X1 U1888 ( .IN1(\ram[67][5] ), .IN2(n566), .IN3(n495), .IN4(n216), .Q(
        n3537) );
  AO22X1 U1889 ( .IN1(\ram[67][6] ), .IN2(n566), .IN3(n495), .IN4(n249), .Q(
        n3538) );
  AO22X1 U1890 ( .IN1(\ram[67][7] ), .IN2(n566), .IN3(n495), .IN4(n282), .Q(
        n3539) );
  AO22X1 U1893 ( .IN1(\ram[66][0] ), .IN2(n569), .IN3(n4136), .IN4(n51), .Q(
        n3540) );
  AO22X1 U1894 ( .IN1(\ram[66][1] ), .IN2(n569), .IN3(n4136), .IN4(n84), .Q(
        n3541) );
  AO22X1 U1895 ( .IN1(\ram[66][2] ), .IN2(n569), .IN3(n4136), .IN4(n117), .Q(
        n3542) );
  AO22X1 U1896 ( .IN1(\ram[66][3] ), .IN2(n569), .IN3(n4136), .IN4(n150), .Q(
        n3543) );
  AO22X1 U1897 ( .IN1(\ram[66][4] ), .IN2(n569), .IN3(n4136), .IN4(n183), .Q(
        n3544) );
  AO22X1 U1898 ( .IN1(\ram[66][5] ), .IN2(n569), .IN3(n4136), .IN4(n216), .Q(
        n3545) );
  AO22X1 U1899 ( .IN1(\ram[66][6] ), .IN2(n569), .IN3(n4136), .IN4(n249), .Q(
        n3546) );
  AO22X1 U1900 ( .IN1(\ram[66][7] ), .IN2(n569), .IN3(n4136), .IN4(n282), .Q(
        n3547) );
  AO22X1 U1903 ( .IN1(\ram[65][0] ), .IN2(n572), .IN3(n591), .IN4(n51), .Q(
        n3548) );
  AO22X1 U1904 ( .IN1(\ram[65][1] ), .IN2(n572), .IN3(n591), .IN4(n84), .Q(
        n3549) );
  AO22X1 U1905 ( .IN1(\ram[65][2] ), .IN2(n572), .IN3(n591), .IN4(n117), .Q(
        n3550) );
  AO22X1 U1906 ( .IN1(\ram[65][3] ), .IN2(n572), .IN3(n591), .IN4(n150), .Q(
        n3551) );
  AO22X1 U1907 ( .IN1(\ram[65][4] ), .IN2(n572), .IN3(n591), .IN4(n183), .Q(
        n3552) );
  AO22X1 U1908 ( .IN1(\ram[65][5] ), .IN2(n572), .IN3(n591), .IN4(n216), .Q(
        n3553) );
  AO22X1 U1909 ( .IN1(\ram[65][6] ), .IN2(n572), .IN3(n591), .IN4(n249), .Q(
        n3554) );
  AO22X1 U1910 ( .IN1(\ram[65][7] ), .IN2(n572), .IN3(n591), .IN4(n282), .Q(
        n3555) );
  AO22X1 U1913 ( .IN1(\ram[64][0] ), .IN2(n575), .IN3(n4125), .IN4(n51), .Q(
        n3556) );
  AO22X1 U1914 ( .IN1(\ram[64][1] ), .IN2(n575), .IN3(n4125), .IN4(n84), .Q(
        n3557) );
  AO22X1 U1915 ( .IN1(\ram[64][2] ), .IN2(n575), .IN3(n4125), .IN4(n117), .Q(
        n3558) );
  AO22X1 U1916 ( .IN1(\ram[64][3] ), .IN2(n575), .IN3(n4125), .IN4(n150), .Q(
        n3559) );
  AO22X1 U1917 ( .IN1(\ram[64][4] ), .IN2(n575), .IN3(n4125), .IN4(n183), .Q(
        n3560) );
  AO22X1 U1918 ( .IN1(\ram[64][5] ), .IN2(n575), .IN3(n4125), .IN4(n216), .Q(
        n3561) );
  AO22X1 U1919 ( .IN1(\ram[64][6] ), .IN2(n575), .IN3(n4125), .IN4(n249), .Q(
        n3562) );
  AO22X1 U1920 ( .IN1(\ram[64][7] ), .IN2(n575), .IN3(n4125), .IN4(n282), .Q(
        n3563) );
  AO22X1 U1923 ( .IN1(\ram[63][0] ), .IN2(n578), .IN3(n366), .IN4(n51), .Q(
        n3564) );
  AO22X1 U1924 ( .IN1(\ram[63][1] ), .IN2(n578), .IN3(n366), .IN4(n84), .Q(
        n3565) );
  AO22X1 U1925 ( .IN1(\ram[63][2] ), .IN2(n578), .IN3(n366), .IN4(n117), .Q(
        n3566) );
  AO22X1 U1926 ( .IN1(\ram[63][3] ), .IN2(n578), .IN3(n366), .IN4(n150), .Q(
        n3567) );
  AO22X1 U1927 ( .IN1(\ram[63][4] ), .IN2(n578), .IN3(n366), .IN4(n183), .Q(
        n3568) );
  AO22X1 U1928 ( .IN1(\ram[63][5] ), .IN2(n578), .IN3(n366), .IN4(n216), .Q(
        n3569) );
  AO22X1 U1929 ( .IN1(\ram[63][6] ), .IN2(n578), .IN3(n366), .IN4(n249), .Q(
        n3570) );
  AO22X1 U1930 ( .IN1(\ram[63][7] ), .IN2(n578), .IN3(n366), .IN4(n282), .Q(
        n3571) );
  AO22X1 U1933 ( .IN1(\ram[62][0] ), .IN2(n581), .IN3(n4096), .IN4(n51), .Q(
        n3572) );
  AO22X1 U1934 ( .IN1(\ram[62][1] ), .IN2(n581), .IN3(n4096), .IN4(n84), .Q(
        n3573) );
  AO22X1 U1935 ( .IN1(\ram[62][2] ), .IN2(n581), .IN3(n4096), .IN4(n117), .Q(
        n3574) );
  AO22X1 U1936 ( .IN1(\ram[62][3] ), .IN2(n581), .IN3(n4096), .IN4(n150), .Q(
        n3575) );
  AO22X1 U1937 ( .IN1(\ram[62][4] ), .IN2(n581), .IN3(n4096), .IN4(n183), .Q(
        n3576) );
  AO22X1 U1938 ( .IN1(\ram[62][5] ), .IN2(n581), .IN3(n4096), .IN4(n216), .Q(
        n3577) );
  AO22X1 U1939 ( .IN1(\ram[62][6] ), .IN2(n581), .IN3(n4096), .IN4(n249), .Q(
        n3578) );
  AO22X1 U1940 ( .IN1(\ram[62][7] ), .IN2(n581), .IN3(n4096), .IN4(n282), .Q(
        n3579) );
  AO22X1 U1943 ( .IN1(\ram[61][0] ), .IN2(n584), .IN3(n471), .IN4(n51), .Q(
        n3580) );
  AO22X1 U1944 ( .IN1(\ram[61][1] ), .IN2(n584), .IN3(n471), .IN4(n84), .Q(
        n3581) );
  AO22X1 U1945 ( .IN1(\ram[61][2] ), .IN2(n584), .IN3(n471), .IN4(n117), .Q(
        n3582) );
  AO22X1 U1946 ( .IN1(\ram[61][3] ), .IN2(n584), .IN3(n471), .IN4(n150), .Q(
        n3583) );
  AO22X1 U1947 ( .IN1(\ram[61][4] ), .IN2(n584), .IN3(n471), .IN4(n183), .Q(
        n3584) );
  AO22X1 U1948 ( .IN1(\ram[61][5] ), .IN2(n584), .IN3(n471), .IN4(n216), .Q(
        n3585) );
  AO22X1 U1949 ( .IN1(\ram[61][6] ), .IN2(n584), .IN3(n471), .IN4(n249), .Q(
        n3586) );
  AO22X1 U1950 ( .IN1(\ram[61][7] ), .IN2(n584), .IN3(n471), .IN4(n282), .Q(
        n3587) );
  AO22X1 U1953 ( .IN1(\ram[60][0] ), .IN2(n587), .IN3(n753), .IN4(n51), .Q(
        n3588) );
  AO22X1 U1954 ( .IN1(\ram[60][1] ), .IN2(n587), .IN3(n753), .IN4(n84), .Q(
        n3589) );
  AO22X1 U1955 ( .IN1(\ram[60][2] ), .IN2(n587), .IN3(n753), .IN4(n117), .Q(
        n3590) );
  AO22X1 U1956 ( .IN1(\ram[60][3] ), .IN2(n587), .IN3(n753), .IN4(n150), .Q(
        n3591) );
  AO22X1 U1957 ( .IN1(\ram[60][4] ), .IN2(n587), .IN3(n753), .IN4(n183), .Q(
        n3592) );
  AO22X1 U1958 ( .IN1(\ram[60][5] ), .IN2(n587), .IN3(n753), .IN4(n216), .Q(
        n3593) );
  AO22X1 U1959 ( .IN1(\ram[60][6] ), .IN2(n587), .IN3(n753), .IN4(n249), .Q(
        n3594) );
  AO22X1 U1960 ( .IN1(\ram[60][7] ), .IN2(n587), .IN3(n753), .IN4(n282), .Q(
        n3595) );
  AO22X1 U1963 ( .IN1(\ram[59][0] ), .IN2(n590), .IN3(n318), .IN4(n48), .Q(
        n3596) );
  AO22X1 U1964 ( .IN1(\ram[59][1] ), .IN2(n590), .IN3(n318), .IN4(n81), .Q(
        n3597) );
  AO22X1 U1965 ( .IN1(\ram[59][2] ), .IN2(n590), .IN3(n318), .IN4(n114), .Q(
        n3598) );
  AO22X1 U1966 ( .IN1(\ram[59][3] ), .IN2(n590), .IN3(n318), .IN4(n147), .Q(
        n3599) );
  AO22X1 U1967 ( .IN1(\ram[59][4] ), .IN2(n590), .IN3(n318), .IN4(n180), .Q(
        n3600) );
  AO22X1 U1968 ( .IN1(\ram[59][5] ), .IN2(n590), .IN3(n318), .IN4(n213), .Q(
        n3601) );
  AO22X1 U1969 ( .IN1(\ram[59][6] ), .IN2(n590), .IN3(n318), .IN4(n246), .Q(
        n3602) );
  AO22X1 U1970 ( .IN1(\ram[59][7] ), .IN2(n590), .IN3(n318), .IN4(n279), .Q(
        n3603) );
  AO22X1 U1973 ( .IN1(\ram[58][0] ), .IN2(n593), .IN3(n4078), .IN4(n48), .Q(
        n3604) );
  AO22X1 U1974 ( .IN1(\ram[58][1] ), .IN2(n593), .IN3(n4078), .IN4(n81), .Q(
        n3605) );
  AO22X1 U1975 ( .IN1(\ram[58][2] ), .IN2(n593), .IN3(n4078), .IN4(n114), .Q(
        n3606) );
  AO22X1 U1976 ( .IN1(\ram[58][3] ), .IN2(n593), .IN3(n4078), .IN4(n147), .Q(
        n3607) );
  AO22X1 U1977 ( .IN1(\ram[58][4] ), .IN2(n593), .IN3(n4078), .IN4(n180), .Q(
        n3608) );
  AO22X1 U1978 ( .IN1(\ram[58][5] ), .IN2(n593), .IN3(n4078), .IN4(n213), .Q(
        n3609) );
  AO22X1 U1979 ( .IN1(\ram[58][6] ), .IN2(n593), .IN3(n4078), .IN4(n246), .Q(
        n3610) );
  AO22X1 U1980 ( .IN1(\ram[58][7] ), .IN2(n593), .IN3(n4078), .IN4(n279), .Q(
        n3611) );
  AO22X1 U1983 ( .IN1(\ram[57][0] ), .IN2(n596), .IN3(n417), .IN4(n48), .Q(
        n3612) );
  AO22X1 U1984 ( .IN1(\ram[57][1] ), .IN2(n596), .IN3(n417), .IN4(n81), .Q(
        n3613) );
  AO22X1 U1985 ( .IN1(\ram[57][2] ), .IN2(n596), .IN3(n417), .IN4(n114), .Q(
        n3614) );
  AO22X1 U1986 ( .IN1(\ram[57][3] ), .IN2(n596), .IN3(n417), .IN4(n147), .Q(
        n3615) );
  AO22X1 U1987 ( .IN1(\ram[57][4] ), .IN2(n596), .IN3(n417), .IN4(n180), .Q(
        n3616) );
  AO22X1 U1988 ( .IN1(\ram[57][5] ), .IN2(n596), .IN3(n417), .IN4(n213), .Q(
        n3617) );
  AO22X1 U1989 ( .IN1(\ram[57][6] ), .IN2(n596), .IN3(n417), .IN4(n246), .Q(
        n3618) );
  AO22X1 U1990 ( .IN1(\ram[57][7] ), .IN2(n596), .IN3(n417), .IN4(n279), .Q(
        n3619) );
  AO22X1 U1993 ( .IN1(\ram[56][0] ), .IN2(n599), .IN3(n705), .IN4(n48), .Q(
        n3620) );
  AO22X1 U1994 ( .IN1(\ram[56][1] ), .IN2(n599), .IN3(n705), .IN4(n81), .Q(
        n3621) );
  AO22X1 U1995 ( .IN1(\ram[56][2] ), .IN2(n599), .IN3(n705), .IN4(n114), .Q(
        n3622) );
  AO22X1 U1996 ( .IN1(\ram[56][3] ), .IN2(n599), .IN3(n705), .IN4(n147), .Q(
        n3623) );
  AO22X1 U1997 ( .IN1(\ram[56][4] ), .IN2(n599), .IN3(n705), .IN4(n180), .Q(
        n3624) );
  AO22X1 U1998 ( .IN1(\ram[56][5] ), .IN2(n599), .IN3(n705), .IN4(n213), .Q(
        n3625) );
  AO22X1 U1999 ( .IN1(\ram[56][6] ), .IN2(n599), .IN3(n705), .IN4(n246), .Q(
        n3626) );
  AO22X1 U2000 ( .IN1(\ram[56][7] ), .IN2(n599), .IN3(n705), .IN4(n279), .Q(
        n3627) );
  AO22X1 U2003 ( .IN1(\ram[55][0] ), .IN2(n602), .IN3(n558), .IN4(n48), .Q(
        n3628) );
  AO22X1 U2004 ( .IN1(\ram[55][1] ), .IN2(n602), .IN3(n558), .IN4(n81), .Q(
        n3629) );
  AO22X1 U2005 ( .IN1(\ram[55][2] ), .IN2(n602), .IN3(n558), .IN4(n114), .Q(
        n3630) );
  AO22X1 U2006 ( .IN1(\ram[55][3] ), .IN2(n602), .IN3(n558), .IN4(n147), .Q(
        n3631) );
  AO22X1 U2007 ( .IN1(\ram[55][4] ), .IN2(n602), .IN3(n558), .IN4(n180), .Q(
        n3632) );
  AO22X1 U2008 ( .IN1(\ram[55][5] ), .IN2(n602), .IN3(n558), .IN4(n213), .Q(
        n3633) );
  AO22X1 U2009 ( .IN1(\ram[55][6] ), .IN2(n602), .IN3(n558), .IN4(n246), .Q(
        n3634) );
  AO22X1 U2010 ( .IN1(\ram[55][7] ), .IN2(n602), .IN3(n558), .IN4(n279), .Q(
        n3635) );
  AO22X1 U2013 ( .IN1(\ram[54][0] ), .IN2(n605), .IN3(n4157), .IN4(n48), .Q(
        n3636) );
  AO22X1 U2014 ( .IN1(\ram[54][1] ), .IN2(n605), .IN3(n4157), .IN4(n81), .Q(
        n3637) );
  AO22X1 U2015 ( .IN1(\ram[54][2] ), .IN2(n605), .IN3(n4157), .IN4(n114), .Q(
        n3638) );
  AO22X1 U2016 ( .IN1(\ram[54][3] ), .IN2(n605), .IN3(n4157), .IN4(n147), .Q(
        n3639) );
  AO22X1 U2017 ( .IN1(\ram[54][4] ), .IN2(n605), .IN3(n4157), .IN4(n180), .Q(
        n3640) );
  AO22X1 U2018 ( .IN1(\ram[54][5] ), .IN2(n605), .IN3(n4157), .IN4(n213), .Q(
        n3641) );
  AO22X1 U2019 ( .IN1(\ram[54][6] ), .IN2(n605), .IN3(n4157), .IN4(n246), .Q(
        n3642) );
  AO22X1 U2020 ( .IN1(\ram[54][7] ), .IN2(n605), .IN3(n4157), .IN4(n279), .Q(
        n3643) );
  AO22X1 U2023 ( .IN1(\ram[53][0] ), .IN2(n608), .IN3(n654), .IN4(n48), .Q(
        n3644) );
  AO22X1 U2024 ( .IN1(\ram[53][1] ), .IN2(n608), .IN3(n654), .IN4(n81), .Q(
        n3645) );
  AO22X1 U2025 ( .IN1(\ram[53][2] ), .IN2(n608), .IN3(n654), .IN4(n114), .Q(
        n3646) );
  AO22X1 U2026 ( .IN1(\ram[53][3] ), .IN2(n608), .IN3(n654), .IN4(n147), .Q(
        n3647) );
  AO22X1 U2027 ( .IN1(\ram[53][4] ), .IN2(n608), .IN3(n654), .IN4(n180), .Q(
        n3648) );
  AO22X1 U2028 ( .IN1(\ram[53][5] ), .IN2(n608), .IN3(n654), .IN4(n213), .Q(
        n3649) );
  AO22X1 U2029 ( .IN1(\ram[53][6] ), .IN2(n608), .IN3(n654), .IN4(n246), .Q(
        n3650) );
  AO22X1 U2030 ( .IN1(\ram[53][7] ), .IN2(n608), .IN3(n654), .IN4(n279), .Q(
        n3651) );
  AO22X1 U2033 ( .IN1(\ram[52][0] ), .IN2(n611), .IN3(n4109), .IN4(n48), .Q(
        n3652) );
  AO22X1 U2034 ( .IN1(\ram[52][1] ), .IN2(n611), .IN3(n4109), .IN4(n81), .Q(
        n3653) );
  AO22X1 U2035 ( .IN1(\ram[52][2] ), .IN2(n611), .IN3(n4109), .IN4(n114), .Q(
        n3654) );
  AO22X1 U2036 ( .IN1(\ram[52][3] ), .IN2(n611), .IN3(n4109), .IN4(n147), .Q(
        n3655) );
  AO22X1 U2037 ( .IN1(\ram[52][4] ), .IN2(n611), .IN3(n4109), .IN4(n180), .Q(
        n3656) );
  AO22X1 U2038 ( .IN1(\ram[52][5] ), .IN2(n611), .IN3(n4109), .IN4(n213), .Q(
        n3657) );
  AO22X1 U2039 ( .IN1(\ram[52][6] ), .IN2(n611), .IN3(n4109), .IN4(n246), .Q(
        n3658) );
  AO22X1 U2040 ( .IN1(\ram[52][7] ), .IN2(n611), .IN3(n4109), .IN4(n279), .Q(
        n3659) );
  AO22X1 U2043 ( .IN1(\ram[51][0] ), .IN2(n614), .IN3(n510), .IN4(n48), .Q(
        n3660) );
  AO22X1 U2044 ( .IN1(\ram[51][1] ), .IN2(n614), .IN3(n510), .IN4(n81), .Q(
        n3661) );
  AO22X1 U2045 ( .IN1(\ram[51][2] ), .IN2(n614), .IN3(n510), .IN4(n114), .Q(
        n3662) );
  AO22X1 U2046 ( .IN1(\ram[51][3] ), .IN2(n614), .IN3(n510), .IN4(n147), .Q(
        n3663) );
  AO22X1 U2047 ( .IN1(\ram[51][4] ), .IN2(n614), .IN3(n510), .IN4(n180), .Q(
        n3664) );
  AO22X1 U2048 ( .IN1(\ram[51][5] ), .IN2(n614), .IN3(n510), .IN4(n213), .Q(
        n3665) );
  AO22X1 U2049 ( .IN1(\ram[51][6] ), .IN2(n614), .IN3(n510), .IN4(n246), .Q(
        n3666) );
  AO22X1 U2050 ( .IN1(\ram[51][7] ), .IN2(n614), .IN3(n510), .IN4(n279), .Q(
        n3667) );
  AO22X1 U2053 ( .IN1(\ram[50][0] ), .IN2(n617), .IN3(n4141), .IN4(n48), .Q(
        n3668) );
  AO22X1 U2054 ( .IN1(\ram[50][1] ), .IN2(n617), .IN3(n4141), .IN4(n81), .Q(
        n3669) );
  AO22X1 U2055 ( .IN1(\ram[50][2] ), .IN2(n617), .IN3(n4141), .IN4(n114), .Q(
        n3670) );
  AO22X1 U2056 ( .IN1(\ram[50][3] ), .IN2(n617), .IN3(n4141), .IN4(n147), .Q(
        n3671) );
  AO22X1 U2057 ( .IN1(\ram[50][4] ), .IN2(n617), .IN3(n4141), .IN4(n180), .Q(
        n3672) );
  AO22X1 U2058 ( .IN1(\ram[50][5] ), .IN2(n617), .IN3(n4141), .IN4(n213), .Q(
        n3673) );
  AO22X1 U2059 ( .IN1(\ram[50][6] ), .IN2(n617), .IN3(n4141), .IN4(n246), .Q(
        n3674) );
  AO22X1 U2060 ( .IN1(\ram[50][7] ), .IN2(n617), .IN3(n4141), .IN4(n279), .Q(
        n3675) );
  AO22X1 U2063 ( .IN1(\ram[49][0] ), .IN2(n620), .IN3(n606), .IN4(n48), .Q(
        n3676) );
  AO22X1 U2064 ( .IN1(\ram[49][1] ), .IN2(n620), .IN3(n606), .IN4(n81), .Q(
        n3677) );
  AO22X1 U2065 ( .IN1(\ram[49][2] ), .IN2(n620), .IN3(n606), .IN4(n114), .Q(
        n3678) );
  AO22X1 U2066 ( .IN1(\ram[49][3] ), .IN2(n620), .IN3(n606), .IN4(n147), .Q(
        n3679) );
  AO22X1 U2067 ( .IN1(\ram[49][4] ), .IN2(n620), .IN3(n606), .IN4(n180), .Q(
        n3680) );
  AO22X1 U2068 ( .IN1(\ram[49][5] ), .IN2(n620), .IN3(n606), .IN4(n213), .Q(
        n3681) );
  AO22X1 U2069 ( .IN1(\ram[49][6] ), .IN2(n620), .IN3(n606), .IN4(n246), .Q(
        n3682) );
  AO22X1 U2070 ( .IN1(\ram[49][7] ), .IN2(n620), .IN3(n606), .IN4(n279), .Q(
        n3683) );
  AO22X1 U2073 ( .IN1(\ram[48][0] ), .IN2(n623), .IN3(n4126), .IN4(n48), .Q(
        n3684) );
  AO22X1 U2074 ( .IN1(\ram[48][1] ), .IN2(n623), .IN3(n4126), .IN4(n81), .Q(
        n3685) );
  AO22X1 U2075 ( .IN1(\ram[48][2] ), .IN2(n623), .IN3(n4126), .IN4(n114), .Q(
        n3686) );
  AO22X1 U2076 ( .IN1(\ram[48][3] ), .IN2(n623), .IN3(n4126), .IN4(n147), .Q(
        n3687) );
  AO22X1 U2077 ( .IN1(\ram[48][4] ), .IN2(n623), .IN3(n4126), .IN4(n180), .Q(
        n3688) );
  AO22X1 U2078 ( .IN1(\ram[48][5] ), .IN2(n623), .IN3(n4126), .IN4(n213), .Q(
        n3689) );
  AO22X1 U2079 ( .IN1(\ram[48][6] ), .IN2(n623), .IN3(n4126), .IN4(n246), .Q(
        n3690) );
  AO22X1 U2080 ( .IN1(\ram[48][7] ), .IN2(n623), .IN3(n4126), .IN4(n279), .Q(
        n3691) );
  AO22X1 U2083 ( .IN1(\ram[47][0] ), .IN2(n626), .IN3(n369), .IN4(n45), .Q(
        n3692) );
  AO22X1 U2084 ( .IN1(\ram[47][1] ), .IN2(n626), .IN3(n369), .IN4(n78), .Q(
        n3693) );
  AO22X1 U2085 ( .IN1(\ram[47][2] ), .IN2(n626), .IN3(n369), .IN4(n111), .Q(
        n3694) );
  AO22X1 U2086 ( .IN1(\ram[47][3] ), .IN2(n626), .IN3(n369), .IN4(n144), .Q(
        n3695) );
  AO22X1 U2087 ( .IN1(\ram[47][4] ), .IN2(n626), .IN3(n369), .IN4(n177), .Q(
        n3696) );
  AO22X1 U2088 ( .IN1(\ram[47][5] ), .IN2(n626), .IN3(n369), .IN4(n210), .Q(
        n3697) );
  AO22X1 U2089 ( .IN1(\ram[47][6] ), .IN2(n626), .IN3(n369), .IN4(n243), .Q(
        n3698) );
  AO22X1 U2090 ( .IN1(\ram[47][7] ), .IN2(n626), .IN3(n369), .IN4(n276), .Q(
        n3699) );
  AO22X1 U2093 ( .IN1(\ram[46][0] ), .IN2(n629), .IN3(n4097), .IN4(n45), .Q(
        n3700) );
  AO22X1 U2094 ( .IN1(\ram[46][1] ), .IN2(n629), .IN3(n4097), .IN4(n78), .Q(
        n3701) );
  AO22X1 U2095 ( .IN1(\ram[46][2] ), .IN2(n629), .IN3(n4097), .IN4(n111), .Q(
        n3702) );
  AO22X1 U2096 ( .IN1(\ram[46][3] ), .IN2(n629), .IN3(n4097), .IN4(n144), .Q(
        n3703) );
  AO22X1 U2097 ( .IN1(\ram[46][4] ), .IN2(n629), .IN3(n4097), .IN4(n177), .Q(
        n3704) );
  AO22X1 U2098 ( .IN1(\ram[46][5] ), .IN2(n629), .IN3(n4097), .IN4(n210), .Q(
        n3705) );
  AO22X1 U2099 ( .IN1(\ram[46][6] ), .IN2(n629), .IN3(n4097), .IN4(n243), .Q(
        n3706) );
  AO22X1 U2100 ( .IN1(\ram[46][7] ), .IN2(n629), .IN3(n4097), .IN4(n276), .Q(
        n3707) );
  AO22X1 U2103 ( .IN1(\ram[45][0] ), .IN2(n632), .IN3(n474), .IN4(n45), .Q(
        n3708) );
  AO22X1 U2104 ( .IN1(\ram[45][1] ), .IN2(n632), .IN3(n474), .IN4(n78), .Q(
        n3709) );
  AO22X1 U2105 ( .IN1(\ram[45][2] ), .IN2(n632), .IN3(n474), .IN4(n111), .Q(
        n3710) );
  AO22X1 U2106 ( .IN1(\ram[45][3] ), .IN2(n632), .IN3(n474), .IN4(n144), .Q(
        n3711) );
  AO22X1 U2107 ( .IN1(\ram[45][4] ), .IN2(n632), .IN3(n474), .IN4(n177), .Q(
        n3712) );
  AO22X1 U2108 ( .IN1(\ram[45][5] ), .IN2(n632), .IN3(n474), .IN4(n210), .Q(
        n3713) );
  AO22X1 U2109 ( .IN1(\ram[45][6] ), .IN2(n632), .IN3(n474), .IN4(n243), .Q(
        n3714) );
  AO22X1 U2110 ( .IN1(\ram[45][7] ), .IN2(n632), .IN3(n474), .IN4(n276), .Q(
        n3715) );
  AO22X1 U2113 ( .IN1(\ram[44][0] ), .IN2(n635), .IN3(n756), .IN4(n45), .Q(
        n3716) );
  AO22X1 U2114 ( .IN1(\ram[44][1] ), .IN2(n635), .IN3(n756), .IN4(n78), .Q(
        n3717) );
  AO22X1 U2115 ( .IN1(\ram[44][2] ), .IN2(n635), .IN3(n756), .IN4(n111), .Q(
        n3718) );
  AO22X1 U2116 ( .IN1(\ram[44][3] ), .IN2(n635), .IN3(n756), .IN4(n144), .Q(
        n3719) );
  AO22X1 U2117 ( .IN1(\ram[44][4] ), .IN2(n635), .IN3(n756), .IN4(n177), .Q(
        n3720) );
  AO22X1 U2118 ( .IN1(\ram[44][5] ), .IN2(n635), .IN3(n756), .IN4(n210), .Q(
        n3721) );
  AO22X1 U2119 ( .IN1(\ram[44][6] ), .IN2(n635), .IN3(n756), .IN4(n243), .Q(
        n3722) );
  AO22X1 U2120 ( .IN1(\ram[44][7] ), .IN2(n635), .IN3(n756), .IN4(n276), .Q(
        n3723) );
  AO22X1 U2123 ( .IN1(\ram[43][0] ), .IN2(n638), .IN3(n321), .IN4(n45), .Q(
        n3724) );
  AO22X1 U2124 ( .IN1(\ram[43][1] ), .IN2(n638), .IN3(n321), .IN4(n78), .Q(
        n3725) );
  AO22X1 U2125 ( .IN1(\ram[43][2] ), .IN2(n638), .IN3(n321), .IN4(n111), .Q(
        n3726) );
  AO22X1 U2126 ( .IN1(\ram[43][3] ), .IN2(n638), .IN3(n321), .IN4(n144), .Q(
        n3727) );
  AO22X1 U2127 ( .IN1(\ram[43][4] ), .IN2(n638), .IN3(n321), .IN4(n177), .Q(
        n3728) );
  AO22X1 U2128 ( .IN1(\ram[43][5] ), .IN2(n638), .IN3(n321), .IN4(n210), .Q(
        n3729) );
  AO22X1 U2129 ( .IN1(\ram[43][6] ), .IN2(n638), .IN3(n321), .IN4(n243), .Q(
        n3730) );
  AO22X1 U2130 ( .IN1(\ram[43][7] ), .IN2(n638), .IN3(n321), .IN4(n276), .Q(
        n3731) );
  AO22X1 U2133 ( .IN1(\ram[42][0] ), .IN2(n641), .IN3(n4079), .IN4(n45), .Q(
        n3732) );
  AO22X1 U2134 ( .IN1(\ram[42][1] ), .IN2(n641), .IN3(n4079), .IN4(n78), .Q(
        n3733) );
  AO22X1 U2135 ( .IN1(\ram[42][2] ), .IN2(n641), .IN3(n4079), .IN4(n111), .Q(
        n3734) );
  AO22X1 U2136 ( .IN1(\ram[42][3] ), .IN2(n641), .IN3(n4079), .IN4(n144), .Q(
        n3735) );
  AO22X1 U2137 ( .IN1(\ram[42][4] ), .IN2(n641), .IN3(n4079), .IN4(n177), .Q(
        n3736) );
  AO22X1 U2138 ( .IN1(\ram[42][5] ), .IN2(n641), .IN3(n4079), .IN4(n210), .Q(
        n3737) );
  AO22X1 U2139 ( .IN1(\ram[42][6] ), .IN2(n641), .IN3(n4079), .IN4(n243), .Q(
        n3738) );
  AO22X1 U2140 ( .IN1(\ram[42][7] ), .IN2(n641), .IN3(n4079), .IN4(n276), .Q(
        n3739) );
  AO22X1 U2143 ( .IN1(\ram[41][0] ), .IN2(n644), .IN3(n420), .IN4(n45), .Q(
        n3740) );
  AO22X1 U2144 ( .IN1(\ram[41][1] ), .IN2(n644), .IN3(n420), .IN4(n78), .Q(
        n3741) );
  AO22X1 U2145 ( .IN1(\ram[41][2] ), .IN2(n644), .IN3(n420), .IN4(n111), .Q(
        n3742) );
  AO22X1 U2146 ( .IN1(\ram[41][3] ), .IN2(n644), .IN3(n420), .IN4(n144), .Q(
        n3743) );
  AO22X1 U2147 ( .IN1(\ram[41][4] ), .IN2(n644), .IN3(n420), .IN4(n177), .Q(
        n3744) );
  AO22X1 U2148 ( .IN1(\ram[41][5] ), .IN2(n644), .IN3(n420), .IN4(n210), .Q(
        n3745) );
  AO22X1 U2149 ( .IN1(\ram[41][6] ), .IN2(n644), .IN3(n420), .IN4(n243), .Q(
        n3746) );
  AO22X1 U2150 ( .IN1(\ram[41][7] ), .IN2(n644), .IN3(n420), .IN4(n276), .Q(
        n3747) );
  AO22X1 U2153 ( .IN1(\ram[40][0] ), .IN2(n647), .IN3(n708), .IN4(n45), .Q(
        n3748) );
  AO22X1 U2154 ( .IN1(\ram[40][1] ), .IN2(n647), .IN3(n708), .IN4(n78), .Q(
        n3749) );
  AO22X1 U2155 ( .IN1(\ram[40][2] ), .IN2(n647), .IN3(n708), .IN4(n111), .Q(
        n3750) );
  AO22X1 U2156 ( .IN1(\ram[40][3] ), .IN2(n647), .IN3(n708), .IN4(n144), .Q(
        n3751) );
  AO22X1 U2157 ( .IN1(\ram[40][4] ), .IN2(n647), .IN3(n708), .IN4(n177), .Q(
        n3752) );
  AO22X1 U2158 ( .IN1(\ram[40][5] ), .IN2(n647), .IN3(n708), .IN4(n210), .Q(
        n3753) );
  AO22X1 U2159 ( .IN1(\ram[40][6] ), .IN2(n647), .IN3(n708), .IN4(n243), .Q(
        n3754) );
  AO22X1 U2160 ( .IN1(\ram[40][7] ), .IN2(n647), .IN3(n708), .IN4(n276), .Q(
        n3755) );
  AO22X1 U2163 ( .IN1(\ram[39][0] ), .IN2(n650), .IN3(n561), .IN4(n45), .Q(
        n3756) );
  AO22X1 U2164 ( .IN1(\ram[39][1] ), .IN2(n650), .IN3(n561), .IN4(n78), .Q(
        n3757) );
  AO22X1 U2165 ( .IN1(\ram[39][2] ), .IN2(n650), .IN3(n561), .IN4(n111), .Q(
        n3758) );
  AO22X1 U2166 ( .IN1(\ram[39][3] ), .IN2(n650), .IN3(n561), .IN4(n144), .Q(
        n3759) );
  AO22X1 U2167 ( .IN1(\ram[39][4] ), .IN2(n650), .IN3(n561), .IN4(n177), .Q(
        n3760) );
  AO22X1 U2168 ( .IN1(\ram[39][5] ), .IN2(n650), .IN3(n561), .IN4(n210), .Q(
        n3761) );
  AO22X1 U2169 ( .IN1(\ram[39][6] ), .IN2(n650), .IN3(n561), .IN4(n243), .Q(
        n3762) );
  AO22X1 U2170 ( .IN1(\ram[39][7] ), .IN2(n650), .IN3(n561), .IN4(n276), .Q(
        n3763) );
  AO22X1 U2173 ( .IN1(\ram[38][0] ), .IN2(n653), .IN3(n4158), .IN4(n45), .Q(
        n3764) );
  AO22X1 U2174 ( .IN1(\ram[38][1] ), .IN2(n653), .IN3(n4158), .IN4(n78), .Q(
        n3765) );
  AO22X1 U2175 ( .IN1(\ram[38][2] ), .IN2(n653), .IN3(n4158), .IN4(n111), .Q(
        n3766) );
  AO22X1 U2176 ( .IN1(\ram[38][3] ), .IN2(n653), .IN3(n4158), .IN4(n144), .Q(
        n3767) );
  AO22X1 U2177 ( .IN1(\ram[38][4] ), .IN2(n653), .IN3(n4158), .IN4(n177), .Q(
        n3768) );
  AO22X1 U2178 ( .IN1(\ram[38][5] ), .IN2(n653), .IN3(n4158), .IN4(n210), .Q(
        n3769) );
  AO22X1 U2179 ( .IN1(\ram[38][6] ), .IN2(n653), .IN3(n4158), .IN4(n243), .Q(
        n3770) );
  AO22X1 U2180 ( .IN1(\ram[38][7] ), .IN2(n653), .IN3(n4158), .IN4(n276), .Q(
        n3771) );
  AO22X1 U2183 ( .IN1(\ram[37][0] ), .IN2(n656), .IN3(n657), .IN4(n45), .Q(
        n3772) );
  AO22X1 U2184 ( .IN1(\ram[37][1] ), .IN2(n656), .IN3(n657), .IN4(n78), .Q(
        n3773) );
  AO22X1 U2185 ( .IN1(\ram[37][2] ), .IN2(n656), .IN3(n657), .IN4(n111), .Q(
        n3774) );
  AO22X1 U2186 ( .IN1(\ram[37][3] ), .IN2(n656), .IN3(n657), .IN4(n144), .Q(
        n3775) );
  AO22X1 U2187 ( .IN1(\ram[37][4] ), .IN2(n656), .IN3(n657), .IN4(n177), .Q(
        n3776) );
  AO22X1 U2188 ( .IN1(\ram[37][5] ), .IN2(n656), .IN3(n657), .IN4(n210), .Q(
        n3777) );
  AO22X1 U2189 ( .IN1(\ram[37][6] ), .IN2(n656), .IN3(n657), .IN4(n243), .Q(
        n3778) );
  AO22X1 U2190 ( .IN1(\ram[37][7] ), .IN2(n656), .IN3(n657), .IN4(n276), .Q(
        n3779) );
  AO22X1 U2193 ( .IN1(\ram[36][0] ), .IN2(n659), .IN3(n4110), .IN4(n45), .Q(
        n3780) );
  AO22X1 U2194 ( .IN1(\ram[36][1] ), .IN2(n659), .IN3(n4110), .IN4(n78), .Q(
        n3781) );
  AO22X1 U2195 ( .IN1(\ram[36][2] ), .IN2(n659), .IN3(n4110), .IN4(n111), .Q(
        n3782) );
  AO22X1 U2196 ( .IN1(\ram[36][3] ), .IN2(n659), .IN3(n4110), .IN4(n144), .Q(
        n3783) );
  AO22X1 U2197 ( .IN1(\ram[36][4] ), .IN2(n659), .IN3(n4110), .IN4(n177), .Q(
        n3784) );
  AO22X1 U2198 ( .IN1(\ram[36][5] ), .IN2(n659), .IN3(n4110), .IN4(n210), .Q(
        n3785) );
  AO22X1 U2199 ( .IN1(\ram[36][6] ), .IN2(n659), .IN3(n4110), .IN4(n243), .Q(
        n3786) );
  AO22X1 U2200 ( .IN1(\ram[36][7] ), .IN2(n659), .IN3(n4110), .IN4(n276), .Q(
        n3787) );
  AO22X1 U2203 ( .IN1(\ram[35][0] ), .IN2(n662), .IN3(n513), .IN4(n42), .Q(
        n3788) );
  AO22X1 U2204 ( .IN1(\ram[35][1] ), .IN2(n662), .IN3(n513), .IN4(n75), .Q(
        n3789) );
  AO22X1 U2205 ( .IN1(\ram[35][2] ), .IN2(n662), .IN3(n513), .IN4(n108), .Q(
        n3790) );
  AO22X1 U2206 ( .IN1(\ram[35][3] ), .IN2(n662), .IN3(n513), .IN4(n141), .Q(
        n3791) );
  AO22X1 U2207 ( .IN1(\ram[35][4] ), .IN2(n662), .IN3(n513), .IN4(n174), .Q(
        n3792) );
  AO22X1 U2208 ( .IN1(\ram[35][5] ), .IN2(n662), .IN3(n513), .IN4(n207), .Q(
        n3793) );
  AO22X1 U2209 ( .IN1(\ram[35][6] ), .IN2(n662), .IN3(n513), .IN4(n240), .Q(
        n3794) );
  AO22X1 U2210 ( .IN1(\ram[35][7] ), .IN2(n662), .IN3(n513), .IN4(n273), .Q(
        n3795) );
  AO22X1 U2213 ( .IN1(\ram[34][0] ), .IN2(n665), .IN3(n4142), .IN4(n42), .Q(
        n3796) );
  AO22X1 U2214 ( .IN1(\ram[34][1] ), .IN2(n665), .IN3(n4142), .IN4(n75), .Q(
        n3797) );
  AO22X1 U2215 ( .IN1(\ram[34][2] ), .IN2(n665), .IN3(n4142), .IN4(n108), .Q(
        n3798) );
  AO22X1 U2216 ( .IN1(\ram[34][3] ), .IN2(n665), .IN3(n4142), .IN4(n141), .Q(
        n3799) );
  AO22X1 U2217 ( .IN1(\ram[34][4] ), .IN2(n665), .IN3(n4142), .IN4(n174), .Q(
        n3800) );
  AO22X1 U2218 ( .IN1(\ram[34][5] ), .IN2(n665), .IN3(n4142), .IN4(n207), .Q(
        n3801) );
  AO22X1 U2219 ( .IN1(\ram[34][6] ), .IN2(n665), .IN3(n4142), .IN4(n240), .Q(
        n3802) );
  AO22X1 U2220 ( .IN1(\ram[34][7] ), .IN2(n665), .IN3(n4142), .IN4(n273), .Q(
        n3803) );
  AO22X1 U2223 ( .IN1(\ram[33][0] ), .IN2(n668), .IN3(n609), .IN4(n42), .Q(
        n3804) );
  AO22X1 U2224 ( .IN1(\ram[33][1] ), .IN2(n668), .IN3(n609), .IN4(n75), .Q(
        n3805) );
  AO22X1 U2225 ( .IN1(\ram[33][2] ), .IN2(n668), .IN3(n609), .IN4(n108), .Q(
        n3806) );
  AO22X1 U2226 ( .IN1(\ram[33][3] ), .IN2(n668), .IN3(n609), .IN4(n141), .Q(
        n3807) );
  AO22X1 U2227 ( .IN1(\ram[33][4] ), .IN2(n668), .IN3(n609), .IN4(n174), .Q(
        n3808) );
  AO22X1 U2228 ( .IN1(\ram[33][5] ), .IN2(n668), .IN3(n609), .IN4(n207), .Q(
        n3809) );
  AO22X1 U2229 ( .IN1(\ram[33][6] ), .IN2(n668), .IN3(n609), .IN4(n240), .Q(
        n3810) );
  AO22X1 U2230 ( .IN1(\ram[33][7] ), .IN2(n668), .IN3(n609), .IN4(n273), .Q(
        n3811) );
  AO22X1 U2233 ( .IN1(\ram[32][0] ), .IN2(n671), .IN3(n4123), .IN4(n42), .Q(
        n3812) );
  AO22X1 U2234 ( .IN1(\ram[32][1] ), .IN2(n671), .IN3(n4123), .IN4(n75), .Q(
        n3813) );
  AO22X1 U2235 ( .IN1(\ram[32][2] ), .IN2(n671), .IN3(n4123), .IN4(n108), .Q(
        n3814) );
  AO22X1 U2236 ( .IN1(\ram[32][3] ), .IN2(n671), .IN3(n4123), .IN4(n141), .Q(
        n3815) );
  AO22X1 U2237 ( .IN1(\ram[32][4] ), .IN2(n671), .IN3(n4123), .IN4(n174), .Q(
        n3816) );
  AO22X1 U2238 ( .IN1(\ram[32][5] ), .IN2(n671), .IN3(n4123), .IN4(n207), .Q(
        n3817) );
  AO22X1 U2239 ( .IN1(\ram[32][6] ), .IN2(n671), .IN3(n4123), .IN4(n240), .Q(
        n3818) );
  AO22X1 U2240 ( .IN1(\ram[32][7] ), .IN2(n671), .IN3(n4123), .IN4(n273), .Q(
        n3819) );
  AO22X1 U2243 ( .IN1(\ram[31][0] ), .IN2(n674), .IN3(n360), .IN4(n42), .Q(
        n3820) );
  AO22X1 U2244 ( .IN1(\ram[31][1] ), .IN2(n674), .IN3(n360), .IN4(n75), .Q(
        n3821) );
  AO22X1 U2245 ( .IN1(\ram[31][2] ), .IN2(n674), .IN3(n360), .IN4(n108), .Q(
        n3822) );
  AO22X1 U2246 ( .IN1(\ram[31][3] ), .IN2(n674), .IN3(n360), .IN4(n141), .Q(
        n3823) );
  AO22X1 U2247 ( .IN1(\ram[31][4] ), .IN2(n674), .IN3(n360), .IN4(n174), .Q(
        n3824) );
  AO22X1 U2248 ( .IN1(\ram[31][5] ), .IN2(n674), .IN3(n360), .IN4(n207), .Q(
        n3825) );
  AO22X1 U2249 ( .IN1(\ram[31][6] ), .IN2(n674), .IN3(n360), .IN4(n240), .Q(
        n3826) );
  AO22X1 U2250 ( .IN1(\ram[31][7] ), .IN2(n674), .IN3(n360), .IN4(n273), .Q(
        n3827) );
  AO22X1 U2253 ( .IN1(\ram[30][0] ), .IN2(n677), .IN3(n4094), .IN4(n42), .Q(
        n3828) );
  AO22X1 U2254 ( .IN1(\ram[30][1] ), .IN2(n677), .IN3(n4094), .IN4(n75), .Q(
        n3829) );
  AO22X1 U2255 ( .IN1(\ram[30][2] ), .IN2(n677), .IN3(n4094), .IN4(n108), .Q(
        n3830) );
  AO22X1 U2256 ( .IN1(\ram[30][3] ), .IN2(n677), .IN3(n4094), .IN4(n141), .Q(
        n3831) );
  AO22X1 U2257 ( .IN1(\ram[30][4] ), .IN2(n677), .IN3(n4094), .IN4(n174), .Q(
        n3832) );
  AO22X1 U2258 ( .IN1(\ram[30][5] ), .IN2(n677), .IN3(n4094), .IN4(n207), .Q(
        n3833) );
  AO22X1 U2259 ( .IN1(\ram[30][6] ), .IN2(n677), .IN3(n4094), .IN4(n240), .Q(
        n3834) );
  AO22X1 U2260 ( .IN1(\ram[30][7] ), .IN2(n677), .IN3(n4094), .IN4(n273), .Q(
        n3835) );
  AO22X1 U2263 ( .IN1(\ram[29][0] ), .IN2(n680), .IN3(n465), .IN4(n42), .Q(
        n3836) );
  AO22X1 U2264 ( .IN1(\ram[29][1] ), .IN2(n680), .IN3(n465), .IN4(n75), .Q(
        n3837) );
  AO22X1 U2265 ( .IN1(\ram[29][2] ), .IN2(n680), .IN3(n465), .IN4(n108), .Q(
        n3838) );
  AO22X1 U2266 ( .IN1(\ram[29][3] ), .IN2(n680), .IN3(n465), .IN4(n141), .Q(
        n3839) );
  AO22X1 U2267 ( .IN1(\ram[29][4] ), .IN2(n680), .IN3(n465), .IN4(n174), .Q(
        n3840) );
  AO22X1 U2268 ( .IN1(\ram[29][5] ), .IN2(n680), .IN3(n465), .IN4(n207), .Q(
        n3841) );
  AO22X1 U2269 ( .IN1(\ram[29][6] ), .IN2(n680), .IN3(n465), .IN4(n240), .Q(
        n3842) );
  AO22X1 U2270 ( .IN1(\ram[29][7] ), .IN2(n680), .IN3(n465), .IN4(n273), .Q(
        n3843) );
  AO22X1 U2273 ( .IN1(\ram[28][0] ), .IN2(n683), .IN3(n747), .IN4(n42), .Q(
        n3844) );
  AO22X1 U2274 ( .IN1(\ram[28][1] ), .IN2(n683), .IN3(n747), .IN4(n75), .Q(
        n3845) );
  AO22X1 U2275 ( .IN1(\ram[28][2] ), .IN2(n683), .IN3(n747), .IN4(n108), .Q(
        n3846) );
  AO22X1 U2276 ( .IN1(\ram[28][3] ), .IN2(n683), .IN3(n747), .IN4(n141), .Q(
        n3847) );
  AO22X1 U2277 ( .IN1(\ram[28][4] ), .IN2(n683), .IN3(n747), .IN4(n174), .Q(
        n3848) );
  AO22X1 U2278 ( .IN1(\ram[28][5] ), .IN2(n683), .IN3(n747), .IN4(n207), .Q(
        n3849) );
  AO22X1 U2279 ( .IN1(\ram[28][6] ), .IN2(n683), .IN3(n747), .IN4(n240), .Q(
        n3850) );
  AO22X1 U2280 ( .IN1(\ram[28][7] ), .IN2(n683), .IN3(n747), .IN4(n273), .Q(
        n3851) );
  AO22X1 U2283 ( .IN1(\ram[27][0] ), .IN2(n686), .IN3(n312), .IN4(n42), .Q(
        n3852) );
  AO22X1 U2284 ( .IN1(\ram[27][1] ), .IN2(n686), .IN3(n312), .IN4(n75), .Q(
        n3853) );
  AO22X1 U2285 ( .IN1(\ram[27][2] ), .IN2(n686), .IN3(n312), .IN4(n108), .Q(
        n3854) );
  AO22X1 U2286 ( .IN1(\ram[27][3] ), .IN2(n686), .IN3(n312), .IN4(n141), .Q(
        n3855) );
  AO22X1 U2287 ( .IN1(\ram[27][4] ), .IN2(n686), .IN3(n312), .IN4(n174), .Q(
        n3856) );
  AO22X1 U2288 ( .IN1(\ram[27][5] ), .IN2(n686), .IN3(n312), .IN4(n207), .Q(
        n3857) );
  AO22X1 U2289 ( .IN1(\ram[27][6] ), .IN2(n686), .IN3(n312), .IN4(n240), .Q(
        n3858) );
  AO22X1 U2290 ( .IN1(\ram[27][7] ), .IN2(n686), .IN3(n312), .IN4(n273), .Q(
        n3859) );
  AO22X1 U2293 ( .IN1(\ram[26][0] ), .IN2(n689), .IN3(n4076), .IN4(n42), .Q(
        n3860) );
  AO22X1 U2294 ( .IN1(\ram[26][1] ), .IN2(n689), .IN3(n4076), .IN4(n75), .Q(
        n3861) );
  AO22X1 U2295 ( .IN1(\ram[26][2] ), .IN2(n689), .IN3(n4076), .IN4(n108), .Q(
        n3862) );
  AO22X1 U2296 ( .IN1(\ram[26][3] ), .IN2(n689), .IN3(n4076), .IN4(n141), .Q(
        n3863) );
  AO22X1 U2297 ( .IN1(\ram[26][4] ), .IN2(n689), .IN3(n4076), .IN4(n174), .Q(
        n3864) );
  AO22X1 U2298 ( .IN1(\ram[26][5] ), .IN2(n689), .IN3(n4076), .IN4(n207), .Q(
        n3865) );
  AO22X1 U2299 ( .IN1(\ram[26][6] ), .IN2(n689), .IN3(n4076), .IN4(n240), .Q(
        n3866) );
  AO22X1 U2300 ( .IN1(\ram[26][7] ), .IN2(n689), .IN3(n4076), .IN4(n273), .Q(
        n3867) );
  AO22X1 U2303 ( .IN1(\ram[25][0] ), .IN2(n692), .IN3(n411), .IN4(n42), .Q(
        n3868) );
  AO22X1 U2304 ( .IN1(\ram[25][1] ), .IN2(n692), .IN3(n411), .IN4(n75), .Q(
        n3869) );
  AO22X1 U2305 ( .IN1(\ram[25][2] ), .IN2(n692), .IN3(n411), .IN4(n108), .Q(
        n3870) );
  AO22X1 U2306 ( .IN1(\ram[25][3] ), .IN2(n692), .IN3(n411), .IN4(n141), .Q(
        n3871) );
  AO22X1 U2307 ( .IN1(\ram[25][4] ), .IN2(n692), .IN3(n411), .IN4(n174), .Q(
        n3872) );
  AO22X1 U2308 ( .IN1(\ram[25][5] ), .IN2(n692), .IN3(n411), .IN4(n207), .Q(
        n3873) );
  AO22X1 U2309 ( .IN1(\ram[25][6] ), .IN2(n692), .IN3(n411), .IN4(n240), .Q(
        n3874) );
  AO22X1 U2310 ( .IN1(\ram[25][7] ), .IN2(n692), .IN3(n411), .IN4(n273), .Q(
        n3875) );
  AO22X1 U2313 ( .IN1(\ram[24][0] ), .IN2(n695), .IN3(n699), .IN4(n42), .Q(
        n3876) );
  AO22X1 U2314 ( .IN1(\ram[24][1] ), .IN2(n695), .IN3(n699), .IN4(n75), .Q(
        n3877) );
  AO22X1 U2315 ( .IN1(\ram[24][2] ), .IN2(n695), .IN3(n699), .IN4(n108), .Q(
        n3878) );
  AO22X1 U2316 ( .IN1(\ram[24][3] ), .IN2(n695), .IN3(n699), .IN4(n141), .Q(
        n3879) );
  AO22X1 U2317 ( .IN1(\ram[24][4] ), .IN2(n695), .IN3(n699), .IN4(n174), .Q(
        n3880) );
  AO22X1 U2318 ( .IN1(\ram[24][5] ), .IN2(n695), .IN3(n699), .IN4(n207), .Q(
        n3881) );
  AO22X1 U2319 ( .IN1(\ram[24][6] ), .IN2(n695), .IN3(n699), .IN4(n240), .Q(
        n3882) );
  AO22X1 U2320 ( .IN1(\ram[24][7] ), .IN2(n695), .IN3(n699), .IN4(n273), .Q(
        n3883) );
  AO22X1 U2323 ( .IN1(\ram[23][0] ), .IN2(n698), .IN3(n552), .IN4(n39), .Q(
        n3884) );
  AO22X1 U2324 ( .IN1(\ram[23][1] ), .IN2(n698), .IN3(n552), .IN4(n72), .Q(
        n3885) );
  AO22X1 U2325 ( .IN1(\ram[23][2] ), .IN2(n698), .IN3(n552), .IN4(n105), .Q(
        n3886) );
  AO22X1 U2326 ( .IN1(\ram[23][3] ), .IN2(n698), .IN3(n552), .IN4(n138), .Q(
        n3887) );
  AO22X1 U2327 ( .IN1(\ram[23][4] ), .IN2(n698), .IN3(n552), .IN4(n171), .Q(
        n3888) );
  AO22X1 U2328 ( .IN1(\ram[23][5] ), .IN2(n698), .IN3(n552), .IN4(n204), .Q(
        n3889) );
  AO22X1 U2329 ( .IN1(\ram[23][6] ), .IN2(n698), .IN3(n552), .IN4(n237), .Q(
        n3890) );
  AO22X1 U2330 ( .IN1(\ram[23][7] ), .IN2(n698), .IN3(n552), .IN4(n270), .Q(
        n3891) );
  AO22X1 U2333 ( .IN1(\ram[22][0] ), .IN2(n701), .IN3(n4155), .IN4(n39), .Q(
        n3892) );
  AO22X1 U2334 ( .IN1(\ram[22][1] ), .IN2(n701), .IN3(n4155), .IN4(n72), .Q(
        n3893) );
  AO22X1 U2335 ( .IN1(\ram[22][2] ), .IN2(n701), .IN3(n4155), .IN4(n105), .Q(
        n3894) );
  AO22X1 U2336 ( .IN1(\ram[22][3] ), .IN2(n701), .IN3(n4155), .IN4(n138), .Q(
        n3895) );
  AO22X1 U2337 ( .IN1(\ram[22][4] ), .IN2(n701), .IN3(n4155), .IN4(n171), .Q(
        n3896) );
  AO22X1 U2338 ( .IN1(\ram[22][5] ), .IN2(n701), .IN3(n4155), .IN4(n204), .Q(
        n3897) );
  AO22X1 U2339 ( .IN1(\ram[22][6] ), .IN2(n701), .IN3(n4155), .IN4(n237), .Q(
        n3898) );
  AO22X1 U2340 ( .IN1(\ram[22][7] ), .IN2(n701), .IN3(n4155), .IN4(n270), .Q(
        n3899) );
  AO22X1 U2343 ( .IN1(\ram[21][0] ), .IN2(n704), .IN3(n648), .IN4(n39), .Q(
        n3900) );
  AO22X1 U2344 ( .IN1(\ram[21][1] ), .IN2(n704), .IN3(n648), .IN4(n72), .Q(
        n3901) );
  AO22X1 U2345 ( .IN1(\ram[21][2] ), .IN2(n704), .IN3(n648), .IN4(n105), .Q(
        n3902) );
  AO22X1 U2346 ( .IN1(\ram[21][3] ), .IN2(n704), .IN3(n648), .IN4(n138), .Q(
        n3903) );
  AO22X1 U2347 ( .IN1(\ram[21][4] ), .IN2(n704), .IN3(n648), .IN4(n171), .Q(
        n3904) );
  AO22X1 U2348 ( .IN1(\ram[21][5] ), .IN2(n704), .IN3(n648), .IN4(n204), .Q(
        n3905) );
  AO22X1 U2349 ( .IN1(\ram[21][6] ), .IN2(n704), .IN3(n648), .IN4(n237), .Q(
        n3906) );
  AO22X1 U2350 ( .IN1(\ram[21][7] ), .IN2(n704), .IN3(n648), .IN4(n270), .Q(
        n3907) );
  AO22X1 U2353 ( .IN1(\ram[20][0] ), .IN2(n707), .IN3(n4107), .IN4(n39), .Q(
        n3908) );
  AO22X1 U2354 ( .IN1(\ram[20][1] ), .IN2(n707), .IN3(n4107), .IN4(n72), .Q(
        n3909) );
  AO22X1 U2355 ( .IN1(\ram[20][2] ), .IN2(n707), .IN3(n4107), .IN4(n105), .Q(
        n3910) );
  AO22X1 U2356 ( .IN1(\ram[20][3] ), .IN2(n707), .IN3(n4107), .IN4(n138), .Q(
        n3911) );
  AO22X1 U2357 ( .IN1(\ram[20][4] ), .IN2(n707), .IN3(n4107), .IN4(n171), .Q(
        n3912) );
  AO22X1 U2358 ( .IN1(\ram[20][5] ), .IN2(n707), .IN3(n4107), .IN4(n204), .Q(
        n3913) );
  AO22X1 U2359 ( .IN1(\ram[20][6] ), .IN2(n707), .IN3(n4107), .IN4(n237), .Q(
        n3914) );
  AO22X1 U2360 ( .IN1(\ram[20][7] ), .IN2(n707), .IN3(n4107), .IN4(n270), .Q(
        n3915) );
  AO22X1 U2363 ( .IN1(\ram[19][0] ), .IN2(n710), .IN3(n504), .IN4(n39), .Q(
        n3916) );
  AO22X1 U2364 ( .IN1(\ram[19][1] ), .IN2(n710), .IN3(n504), .IN4(n72), .Q(
        n3917) );
  AO22X1 U2365 ( .IN1(\ram[19][2] ), .IN2(n710), .IN3(n504), .IN4(n105), .Q(
        n3918) );
  AO22X1 U2366 ( .IN1(\ram[19][3] ), .IN2(n710), .IN3(n504), .IN4(n138), .Q(
        n3919) );
  AO22X1 U2367 ( .IN1(\ram[19][4] ), .IN2(n710), .IN3(n504), .IN4(n171), .Q(
        n3920) );
  AO22X1 U2368 ( .IN1(\ram[19][5] ), .IN2(n710), .IN3(n504), .IN4(n204), .Q(
        n3921) );
  AO22X1 U2369 ( .IN1(\ram[19][6] ), .IN2(n710), .IN3(n504), .IN4(n237), .Q(
        n3922) );
  AO22X1 U2370 ( .IN1(\ram[19][7] ), .IN2(n710), .IN3(n504), .IN4(n270), .Q(
        n3923) );
  AO22X1 U2373 ( .IN1(\ram[18][0] ), .IN2(n713), .IN3(n4139), .IN4(n39), .Q(
        n3924) );
  AO22X1 U2374 ( .IN1(\ram[18][1] ), .IN2(n713), .IN3(n4139), .IN4(n72), .Q(
        n3925) );
  AO22X1 U2375 ( .IN1(\ram[18][2] ), .IN2(n713), .IN3(n4139), .IN4(n105), .Q(
        n3926) );
  AO22X1 U2376 ( .IN1(\ram[18][3] ), .IN2(n713), .IN3(n4139), .IN4(n138), .Q(
        n3927) );
  AO22X1 U2377 ( .IN1(\ram[18][4] ), .IN2(n713), .IN3(n4139), .IN4(n171), .Q(
        n3928) );
  AO22X1 U2378 ( .IN1(\ram[18][5] ), .IN2(n713), .IN3(n4139), .IN4(n204), .Q(
        n3929) );
  AO22X1 U2379 ( .IN1(\ram[18][6] ), .IN2(n713), .IN3(n4139), .IN4(n237), .Q(
        n3930) );
  AO22X1 U2380 ( .IN1(\ram[18][7] ), .IN2(n713), .IN3(n4139), .IN4(n270), .Q(
        n3931) );
  AO22X1 U2383 ( .IN1(\ram[17][0] ), .IN2(n716), .IN3(n600), .IN4(n39), .Q(
        n3932) );
  AO22X1 U2384 ( .IN1(\ram[17][1] ), .IN2(n716), .IN3(n600), .IN4(n72), .Q(
        n3933) );
  AO22X1 U2385 ( .IN1(\ram[17][2] ), .IN2(n716), .IN3(n600), .IN4(n105), .Q(
        n3934) );
  AO22X1 U2386 ( .IN1(\ram[17][3] ), .IN2(n716), .IN3(n600), .IN4(n138), .Q(
        n3935) );
  AO22X1 U2387 ( .IN1(\ram[17][4] ), .IN2(n716), .IN3(n600), .IN4(n171), .Q(
        n3936) );
  AO22X1 U2388 ( .IN1(\ram[17][5] ), .IN2(n716), .IN3(n600), .IN4(n204), .Q(
        n3937) );
  AO22X1 U2389 ( .IN1(\ram[17][6] ), .IN2(n716), .IN3(n600), .IN4(n237), .Q(
        n3938) );
  AO22X1 U2390 ( .IN1(\ram[17][7] ), .IN2(n716), .IN3(n600), .IN4(n270), .Q(
        n3939) );
  AO22X1 U2393 ( .IN1(\ram[16][0] ), .IN2(n719), .IN3(n4124), .IN4(n39), .Q(
        n3940) );
  AO22X1 U2394 ( .IN1(\ram[16][1] ), .IN2(n719), .IN3(n4124), .IN4(n72), .Q(
        n3941) );
  AO22X1 U2395 ( .IN1(\ram[16][2] ), .IN2(n719), .IN3(n4124), .IN4(n105), .Q(
        n3942) );
  AO22X1 U2396 ( .IN1(\ram[16][3] ), .IN2(n719), .IN3(n4124), .IN4(n138), .Q(
        n3943) );
  AO22X1 U2397 ( .IN1(\ram[16][4] ), .IN2(n719), .IN3(n4124), .IN4(n171), .Q(
        n3944) );
  AO22X1 U2398 ( .IN1(\ram[16][5] ), .IN2(n719), .IN3(n4124), .IN4(n204), .Q(
        n3945) );
  AO22X1 U2399 ( .IN1(\ram[16][6] ), .IN2(n719), .IN3(n4124), .IN4(n237), .Q(
        n3946) );
  AO22X1 U2400 ( .IN1(\ram[16][7] ), .IN2(n719), .IN3(n4124), .IN4(n270), .Q(
        n3947) );
  AO22X1 U2403 ( .IN1(\ram[15][0] ), .IN2(n722), .IN3(n363), .IN4(n39), .Q(
        n3948) );
  AO22X1 U2404 ( .IN1(\ram[15][1] ), .IN2(n722), .IN3(n363), .IN4(n72), .Q(
        n3949) );
  AO22X1 U2405 ( .IN1(\ram[15][2] ), .IN2(n722), .IN3(n363), .IN4(n105), .Q(
        n3950) );
  AO22X1 U2406 ( .IN1(\ram[15][3] ), .IN2(n722), .IN3(n363), .IN4(n138), .Q(
        n3951) );
  AO22X1 U2407 ( .IN1(\ram[15][4] ), .IN2(n722), .IN3(n363), .IN4(n171), .Q(
        n3952) );
  AO22X1 U2408 ( .IN1(\ram[15][5] ), .IN2(n722), .IN3(n363), .IN4(n204), .Q(
        n3953) );
  AO22X1 U2409 ( .IN1(\ram[15][6] ), .IN2(n722), .IN3(n363), .IN4(n237), .Q(
        n3954) );
  AO22X1 U2410 ( .IN1(\ram[15][7] ), .IN2(n722), .IN3(n363), .IN4(n270), .Q(
        n3955) );
  AO22X1 U2413 ( .IN1(\ram[14][0] ), .IN2(n725), .IN3(n4095), .IN4(n39), .Q(
        n3956) );
  AO22X1 U2414 ( .IN1(\ram[14][1] ), .IN2(n725), .IN3(n4095), .IN4(n72), .Q(
        n3957) );
  AO22X1 U2415 ( .IN1(\ram[14][2] ), .IN2(n725), .IN3(n4095), .IN4(n105), .Q(
        n3958) );
  AO22X1 U2416 ( .IN1(\ram[14][3] ), .IN2(n725), .IN3(n4095), .IN4(n138), .Q(
        n3959) );
  AO22X1 U2417 ( .IN1(\ram[14][4] ), .IN2(n725), .IN3(n4095), .IN4(n171), .Q(
        n3960) );
  AO22X1 U2418 ( .IN1(\ram[14][5] ), .IN2(n725), .IN3(n4095), .IN4(n204), .Q(
        n3961) );
  AO22X1 U2419 ( .IN1(\ram[14][6] ), .IN2(n725), .IN3(n4095), .IN4(n237), .Q(
        n3962) );
  AO22X1 U2420 ( .IN1(\ram[14][7] ), .IN2(n725), .IN3(n4095), .IN4(n270), .Q(
        n3963) );
  AO22X1 U2423 ( .IN1(\ram[13][0] ), .IN2(n728), .IN3(n468), .IN4(n39), .Q(
        n3964) );
  AO22X1 U2424 ( .IN1(\ram[13][1] ), .IN2(n728), .IN3(n468), .IN4(n72), .Q(
        n3965) );
  AO22X1 U2425 ( .IN1(\ram[13][2] ), .IN2(n728), .IN3(n468), .IN4(n105), .Q(
        n3966) );
  AO22X1 U2426 ( .IN1(\ram[13][3] ), .IN2(n728), .IN3(n468), .IN4(n138), .Q(
        n3967) );
  AO22X1 U2427 ( .IN1(\ram[13][4] ), .IN2(n728), .IN3(n468), .IN4(n171), .Q(
        n3968) );
  AO22X1 U2428 ( .IN1(\ram[13][5] ), .IN2(n728), .IN3(n468), .IN4(n204), .Q(
        n3969) );
  AO22X1 U2429 ( .IN1(\ram[13][6] ), .IN2(n728), .IN3(n468), .IN4(n237), .Q(
        n3970) );
  AO22X1 U2430 ( .IN1(\ram[13][7] ), .IN2(n728), .IN3(n468), .IN4(n270), .Q(
        n3971) );
  AO22X1 U2433 ( .IN1(\ram[12][0] ), .IN2(n731), .IN3(n750), .IN4(n39), .Q(
        n3972) );
  AO22X1 U2434 ( .IN1(\ram[12][1] ), .IN2(n731), .IN3(n750), .IN4(n72), .Q(
        n3973) );
  AO22X1 U2435 ( .IN1(\ram[12][2] ), .IN2(n731), .IN3(n750), .IN4(n105), .Q(
        n3974) );
  AO22X1 U2436 ( .IN1(\ram[12][3] ), .IN2(n731), .IN3(n750), .IN4(n138), .Q(
        n3975) );
  AO22X1 U2437 ( .IN1(\ram[12][4] ), .IN2(n731), .IN3(n750), .IN4(n171), .Q(
        n3976) );
  AO22X1 U2438 ( .IN1(\ram[12][5] ), .IN2(n731), .IN3(n750), .IN4(n204), .Q(
        n3977) );
  AO22X1 U2439 ( .IN1(\ram[12][6] ), .IN2(n731), .IN3(n750), .IN4(n237), .Q(
        n3978) );
  AO22X1 U2440 ( .IN1(\ram[12][7] ), .IN2(n731), .IN3(n750), .IN4(n270), .Q(
        n3979) );
  AO22X1 U2443 ( .IN1(\ram[11][0] ), .IN2(n734), .IN3(n315), .IN4(n36), .Q(
        n3980) );
  AO22X1 U2444 ( .IN1(\ram[11][1] ), .IN2(n734), .IN3(n315), .IN4(n69), .Q(
        n3981) );
  AO22X1 U2445 ( .IN1(\ram[11][2] ), .IN2(n734), .IN3(n315), .IN4(n102), .Q(
        n3982) );
  AO22X1 U2446 ( .IN1(\ram[11][3] ), .IN2(n734), .IN3(n315), .IN4(n135), .Q(
        n3983) );
  AO22X1 U2447 ( .IN1(\ram[11][4] ), .IN2(n734), .IN3(n315), .IN4(n168), .Q(
        n3984) );
  AO22X1 U2448 ( .IN1(\ram[11][5] ), .IN2(n734), .IN3(n315), .IN4(n201), .Q(
        n3985) );
  AO22X1 U2449 ( .IN1(\ram[11][6] ), .IN2(n734), .IN3(n315), .IN4(n234), .Q(
        n3986) );
  AO22X1 U2450 ( .IN1(\ram[11][7] ), .IN2(n734), .IN3(n315), .IN4(n267), .Q(
        n3987) );
  AO22X1 U2453 ( .IN1(\ram[10][0] ), .IN2(n737), .IN3(n4077), .IN4(n36), .Q(
        n3988) );
  AO22X1 U2454 ( .IN1(\ram[10][1] ), .IN2(n737), .IN3(n4077), .IN4(n69), .Q(
        n3989) );
  AO22X1 U2455 ( .IN1(\ram[10][2] ), .IN2(n737), .IN3(n4077), .IN4(n102), .Q(
        n3990) );
  AO22X1 U2456 ( .IN1(\ram[10][3] ), .IN2(n737), .IN3(n4077), .IN4(n135), .Q(
        n3991) );
  AO22X1 U2457 ( .IN1(\ram[10][4] ), .IN2(n737), .IN3(n4077), .IN4(n168), .Q(
        n3992) );
  AO22X1 U2458 ( .IN1(\ram[10][5] ), .IN2(n737), .IN3(n4077), .IN4(n201), .Q(
        n3993) );
  AO22X1 U2459 ( .IN1(\ram[10][6] ), .IN2(n737), .IN3(n4077), .IN4(n234), .Q(
        n3994) );
  AO22X1 U2460 ( .IN1(\ram[10][7] ), .IN2(n737), .IN3(n4077), .IN4(n267), .Q(
        n3995) );
  AO22X1 U2463 ( .IN1(\ram[9][0] ), .IN2(n740), .IN3(n414), .IN4(n36), .Q(
        n3996) );
  AO22X1 U2464 ( .IN1(\ram[9][1] ), .IN2(n740), .IN3(n414), .IN4(n69), .Q(
        n3997) );
  AO22X1 U2465 ( .IN1(\ram[9][2] ), .IN2(n740), .IN3(n414), .IN4(n102), .Q(
        n3998) );
  AO22X1 U2466 ( .IN1(\ram[9][3] ), .IN2(n740), .IN3(n414), .IN4(n135), .Q(
        n3999) );
  AO22X1 U2467 ( .IN1(\ram[9][4] ), .IN2(n740), .IN3(n414), .IN4(n168), .Q(
        n4000) );
  AO22X1 U2468 ( .IN1(\ram[9][5] ), .IN2(n740), .IN3(n414), .IN4(n201), .Q(
        n4001) );
  AO22X1 U2469 ( .IN1(\ram[9][6] ), .IN2(n740), .IN3(n414), .IN4(n234), .Q(
        n4002) );
  AO22X1 U2470 ( .IN1(\ram[9][7] ), .IN2(n740), .IN3(n414), .IN4(n267), .Q(
        n4003) );
  AO22X1 U2473 ( .IN1(\ram[8][0] ), .IN2(n743), .IN3(n702), .IN4(n36), .Q(
        n4004) );
  AO22X1 U2474 ( .IN1(\ram[8][1] ), .IN2(n743), .IN3(n702), .IN4(n69), .Q(
        n4005) );
  AO22X1 U2475 ( .IN1(\ram[8][2] ), .IN2(n743), .IN3(n702), .IN4(n102), .Q(
        n4006) );
  AO22X1 U2476 ( .IN1(\ram[8][3] ), .IN2(n743), .IN3(n702), .IN4(n135), .Q(
        n4007) );
  AO22X1 U2477 ( .IN1(\ram[8][4] ), .IN2(n743), .IN3(n702), .IN4(n168), .Q(
        n4008) );
  AO22X1 U2478 ( .IN1(\ram[8][5] ), .IN2(n743), .IN3(n702), .IN4(n201), .Q(
        n4009) );
  AO22X1 U2479 ( .IN1(\ram[8][6] ), .IN2(n743), .IN3(n702), .IN4(n234), .Q(
        n4010) );
  AO22X1 U2480 ( .IN1(\ram[8][7] ), .IN2(n743), .IN3(n702), .IN4(n267), .Q(
        n4011) );
  AO22X1 U2483 ( .IN1(\ram[7][0] ), .IN2(n746), .IN3(n555), .IN4(n36), .Q(
        n4012) );
  AO22X1 U2484 ( .IN1(\ram[7][1] ), .IN2(n746), .IN3(n555), .IN4(n69), .Q(
        n4013) );
  AO22X1 U2485 ( .IN1(\ram[7][2] ), .IN2(n746), .IN3(n555), .IN4(n102), .Q(
        n4014) );
  AO22X1 U2486 ( .IN1(\ram[7][3] ), .IN2(n746), .IN3(n555), .IN4(n135), .Q(
        n4015) );
  AO22X1 U2487 ( .IN1(\ram[7][4] ), .IN2(n746), .IN3(n555), .IN4(n168), .Q(
        n4016) );
  AO22X1 U2488 ( .IN1(\ram[7][5] ), .IN2(n746), .IN3(n555), .IN4(n201), .Q(
        n4017) );
  AO22X1 U2489 ( .IN1(\ram[7][6] ), .IN2(n746), .IN3(n555), .IN4(n234), .Q(
        n4018) );
  AO22X1 U2490 ( .IN1(\ram[7][7] ), .IN2(n746), .IN3(n555), .IN4(n267), .Q(
        n4019) );
  AO22X1 U2493 ( .IN1(\ram[6][0] ), .IN2(n749), .IN3(n4156), .IN4(n36), .Q(
        n4020) );
  AO22X1 U2494 ( .IN1(\ram[6][1] ), .IN2(n749), .IN3(n4156), .IN4(n69), .Q(
        n4021) );
  AO22X1 U2495 ( .IN1(\ram[6][2] ), .IN2(n749), .IN3(n4156), .IN4(n102), .Q(
        n4022) );
  AO22X1 U2496 ( .IN1(\ram[6][3] ), .IN2(n749), .IN3(n4156), .IN4(n135), .Q(
        n4023) );
  AO22X1 U2497 ( .IN1(\ram[6][4] ), .IN2(n749), .IN3(n4156), .IN4(n168), .Q(
        n4024) );
  AO22X1 U2498 ( .IN1(\ram[6][5] ), .IN2(n749), .IN3(n4156), .IN4(n201), .Q(
        n4025) );
  AO22X1 U2499 ( .IN1(\ram[6][6] ), .IN2(n749), .IN3(n4156), .IN4(n234), .Q(
        n4026) );
  AO22X1 U2500 ( .IN1(\ram[6][7] ), .IN2(n749), .IN3(n4156), .IN4(n267), .Q(
        n4027) );
  AO22X1 U2503 ( .IN1(\ram[5][0] ), .IN2(n752), .IN3(n651), .IN4(n36), .Q(
        n4028) );
  AO22X1 U2504 ( .IN1(\ram[5][1] ), .IN2(n752), .IN3(n651), .IN4(n69), .Q(
        n4029) );
  AO22X1 U2505 ( .IN1(\ram[5][2] ), .IN2(n752), .IN3(n651), .IN4(n102), .Q(
        n4030) );
  AO22X1 U2506 ( .IN1(\ram[5][3] ), .IN2(n752), .IN3(n651), .IN4(n135), .Q(
        n4031) );
  AO22X1 U2507 ( .IN1(\ram[5][4] ), .IN2(n752), .IN3(n651), .IN4(n168), .Q(
        n4032) );
  AO22X1 U2508 ( .IN1(\ram[5][5] ), .IN2(n752), .IN3(n651), .IN4(n201), .Q(
        n4033) );
  AO22X1 U2509 ( .IN1(\ram[5][6] ), .IN2(n752), .IN3(n651), .IN4(n234), .Q(
        n4034) );
  AO22X1 U2510 ( .IN1(\ram[5][7] ), .IN2(n752), .IN3(n651), .IN4(n267), .Q(
        n4035) );
  AO22X1 U2513 ( .IN1(\ram[4][0] ), .IN2(n755), .IN3(n4108), .IN4(n36), .Q(
        n4036) );
  AO22X1 U2514 ( .IN1(\ram[4][1] ), .IN2(n755), .IN3(n4108), .IN4(n69), .Q(
        n4037) );
  AO22X1 U2515 ( .IN1(\ram[4][2] ), .IN2(n755), .IN3(n4108), .IN4(n102), .Q(
        n4038) );
  AO22X1 U2516 ( .IN1(\ram[4][3] ), .IN2(n755), .IN3(n4108), .IN4(n135), .Q(
        n4039) );
  AO22X1 U2517 ( .IN1(\ram[4][4] ), .IN2(n755), .IN3(n4108), .IN4(n168), .Q(
        n4040) );
  AO22X1 U2518 ( .IN1(\ram[4][5] ), .IN2(n755), .IN3(n4108), .IN4(n201), .Q(
        n4041) );
  AO22X1 U2519 ( .IN1(\ram[4][6] ), .IN2(n755), .IN3(n4108), .IN4(n234), .Q(
        n4042) );
  AO22X1 U2520 ( .IN1(\ram[4][7] ), .IN2(n755), .IN3(n4108), .IN4(n267), .Q(
        n4043) );
  AO22X1 U2523 ( .IN1(\ram[3][0] ), .IN2(n758), .IN3(n507), .IN4(n36), .Q(
        n4044) );
  AO22X1 U2524 ( .IN1(\ram[3][1] ), .IN2(n758), .IN3(n507), .IN4(n69), .Q(
        n4045) );
  AO22X1 U2525 ( .IN1(\ram[3][2] ), .IN2(n758), .IN3(n507), .IN4(n102), .Q(
        n4046) );
  AO22X1 U2526 ( .IN1(\ram[3][3] ), .IN2(n758), .IN3(n507), .IN4(n135), .Q(
        n4047) );
  AO22X1 U2527 ( .IN1(\ram[3][4] ), .IN2(n758), .IN3(n507), .IN4(n168), .Q(
        n4048) );
  AO22X1 U2528 ( .IN1(\ram[3][5] ), .IN2(n758), .IN3(n507), .IN4(n201), .Q(
        n4049) );
  AO22X1 U2529 ( .IN1(\ram[3][6] ), .IN2(n758), .IN3(n507), .IN4(n234), .Q(
        n4050) );
  AO22X1 U2530 ( .IN1(\ram[3][7] ), .IN2(n758), .IN3(n507), .IN4(n267), .Q(
        n4051) );
  AO22X1 U2533 ( .IN1(\ram[2][0] ), .IN2(n761), .IN3(n4140), .IN4(n36), .Q(
        n4052) );
  AO22X1 U2534 ( .IN1(\ram[2][1] ), .IN2(n761), .IN3(n4140), .IN4(n69), .Q(
        n4053) );
  AO22X1 U2535 ( .IN1(\ram[2][2] ), .IN2(n761), .IN3(n4140), .IN4(n102), .Q(
        n4054) );
  AO22X1 U2536 ( .IN1(\ram[2][3] ), .IN2(n761), .IN3(n4140), .IN4(n135), .Q(
        n4055) );
  AO22X1 U2537 ( .IN1(\ram[2][4] ), .IN2(n761), .IN3(n4140), .IN4(n168), .Q(
        n4056) );
  AO22X1 U2538 ( .IN1(\ram[2][5] ), .IN2(n761), .IN3(n4140), .IN4(n201), .Q(
        n4057) );
  AO22X1 U2539 ( .IN1(\ram[2][6] ), .IN2(n761), .IN3(n4140), .IN4(n234), .Q(
        n4058) );
  AO22X1 U2540 ( .IN1(\ram[2][7] ), .IN2(n761), .IN3(n4140), .IN4(n267), .Q(
        n4059) );
  AO22X1 U2543 ( .IN1(\ram[1][0] ), .IN2(n764), .IN3(n603), .IN4(n36), .Q(
        n4060) );
  AO22X1 U2544 ( .IN1(\ram[1][1] ), .IN2(n764), .IN3(n603), .IN4(n69), .Q(
        n4061) );
  AO22X1 U2545 ( .IN1(\ram[1][2] ), .IN2(n764), .IN3(n603), .IN4(n102), .Q(
        n4062) );
  AO22X1 U2546 ( .IN1(\ram[1][3] ), .IN2(n764), .IN3(n603), .IN4(n135), .Q(
        n4063) );
  AO22X1 U2547 ( .IN1(\ram[1][4] ), .IN2(n764), .IN3(n603), .IN4(n168), .Q(
        n4064) );
  AO22X1 U2548 ( .IN1(\ram[1][5] ), .IN2(n764), .IN3(n603), .IN4(n201), .Q(
        n4065) );
  AO22X1 U2549 ( .IN1(\ram[1][6] ), .IN2(n764), .IN3(n603), .IN4(n234), .Q(
        n4066) );
  AO22X1 U2550 ( .IN1(\ram[1][7] ), .IN2(n764), .IN3(n603), .IN4(n267), .Q(
        n4067) );
  AO22X1 U2553 ( .IN1(\ram[0][0] ), .IN2(n767), .IN3(n4132), .IN4(n36), .Q(
        n4068) );
  AO22X1 U2554 ( .IN1(\ram[0][1] ), .IN2(n767), .IN3(n4132), .IN4(n69), .Q(
        n4069) );
  AO22X1 U2555 ( .IN1(\ram[0][2] ), .IN2(n767), .IN3(n4132), .IN4(n102), .Q(
        n4070) );
  AO22X1 U2556 ( .IN1(\ram[0][3] ), .IN2(n767), .IN3(n4132), .IN4(n135), .Q(
        n4071) );
  AO22X1 U2557 ( .IN1(\ram[0][4] ), .IN2(n767), .IN3(n4132), .IN4(n168), .Q(
        n4072) );
  AO22X1 U2558 ( .IN1(\ram[0][5] ), .IN2(n767), .IN3(n4132), .IN4(n201), .Q(
        n4073) );
  AO22X1 U2559 ( .IN1(\ram[0][6] ), .IN2(n767), .IN3(n4132), .IN4(n234), .Q(
        n4074) );
  AO22X1 U2560 ( .IN1(\ram[0][7] ), .IN2(n767), .IN3(n4132), .IN4(n267), .Q(
        n4075) );
  AO22X1 U2564 ( .IN1(n771), .IN2(dataout[0]), .IN3(n4174), .IN4(n772), .Q(
        n2020) );
  NAND4X0 U2565 ( .IN1(n773), .IN2(n774), .IN3(n775), .IN4(n776), .QN(n772) );
  NAND4X0 U2567 ( .IN1(n781), .IN2(n782), .IN3(n783), .IN4(n784), .QN(n780) );
  AOI221X1 U2568 ( .IN1(n259), .IN2(\ram[170][0] ), .IN3(n262), .IN4(
        \ram[169][0] ), .IN5(n785), .QN(n784) );
  AO22X1 U2569 ( .IN1(n250), .IN2(\ram[173][0] ), .IN3(n247), .IN4(
        \ram[174][0] ), .Q(n785) );
  AOI221X1 U2570 ( .IN1(n283), .IN2(\ram[162][0] ), .IN3(n286), .IN4(
        \ram[161][0] ), .IN5(n786), .QN(n783) );
  AO22X1 U2571 ( .IN1(n274), .IN2(\ram[165][0] ), .IN3(n271), .IN4(
        \ram[166][0] ), .Q(n786) );
  AOI221X1 U2572 ( .IN1(n211), .IN2(\ram[186][0] ), .IN3(n214), .IN4(
        \ram[185][0] ), .IN5(n787), .QN(n782) );
  AO22X1 U2573 ( .IN1(n196), .IN2(\ram[191][0] ), .IN3(n193), .IN4(
        \ram[192][0] ), .Q(n787) );
  AOI221X1 U2574 ( .IN1(n235), .IN2(\ram[178][0] ), .IN3(n238), .IN4(
        \ram[177][0] ), .IN5(n788), .QN(n781) );
  AO22X1 U2575 ( .IN1(n226), .IN2(\ram[181][0] ), .IN3(n223), .IN4(
        \ram[182][0] ), .Q(n788) );
  NAND4X0 U2576 ( .IN1(n789), .IN2(n790), .IN3(n791), .IN4(n792), .QN(n779) );
  AOI221X1 U2577 ( .IN1(n355), .IN2(\ram[138][0] ), .IN3(n358), .IN4(
        \ram[137][0] ), .IN5(n793), .QN(n792) );
  AO22X1 U2578 ( .IN1(n346), .IN2(\ram[141][0] ), .IN3(n343), .IN4(
        \ram[142][0] ), .Q(n793) );
  AOI221X1 U2579 ( .IN1(n379), .IN2(\ram[130][0] ), .IN3(n382), .IN4(
        \ram[129][0] ), .IN5(n794), .QN(n791) );
  AO22X1 U2580 ( .IN1(n370), .IN2(\ram[133][0] ), .IN3(n367), .IN4(
        \ram[134][0] ), .Q(n794) );
  AOI221X1 U2581 ( .IN1(n307), .IN2(\ram[154][0] ), .IN3(n310), .IN4(
        \ram[153][0] ), .IN5(n795), .QN(n790) );
  AO22X1 U2582 ( .IN1(n298), .IN2(\ram[157][0] ), .IN3(n295), .IN4(
        \ram[158][0] ), .Q(n795) );
  AOI221X1 U2583 ( .IN1(n331), .IN2(\ram[146][0] ), .IN3(n334), .IN4(
        \ram[145][0] ), .IN5(n796), .QN(n789) );
  AO22X1 U2584 ( .IN1(n322), .IN2(\ram[149][0] ), .IN3(n319), .IN4(
        \ram[150][0] ), .Q(n796) );
  NAND4X0 U2585 ( .IN1(n797), .IN2(n798), .IN3(n799), .IN4(n800), .QN(n778) );
  AOI221X1 U2586 ( .IN1(n70), .IN2(\ram[233][0] ), .IN3(n49), .IN4(
        \ram[240][0] ), .IN5(n801), .QN(n800) );
  AO22X1 U2587 ( .IN1(n139), .IN2(\ram[210][0] ), .IN3(n52), .IN4(
        \ram[239][0] ), .Q(n801) );
  AOI221X1 U2588 ( .IN1(n94), .IN2(\ram[225][0] ), .IN3(n79), .IN4(
        \ram[230][0] ), .IN5(n802), .QN(n799) );
  AO22X1 U2589 ( .IN1(n67), .IN2(\ram[234][0] ), .IN3(n82), .IN4(\ram[229][0] ), .Q(n802) );
  AOI221X1 U2590 ( .IN1(n13), .IN2(\ram[252][0] ), .IN3(n16), .IN4(
        \ram[251][0] ), .IN5(n803), .QN(n798) );
  AO22X1 U2591 ( .IN1(n91), .IN2(\ram[226][0] ), .IN3(n3), .IN4(\ram[255][0] ), 
        .Q(n803) );
  AOI221X1 U2592 ( .IN1(n43), .IN2(\ram[242][0] ), .IN3(n46), .IN4(
        \ram[241][0] ), .IN5(n804), .QN(n797) );
  AO22X1 U2593 ( .IN1(n34), .IN2(\ram[245][0] ), .IN3(n31), .IN4(\ram[246][0] ), .Q(n804) );
  NAND4X0 U2594 ( .IN1(n805), .IN2(n806), .IN3(n807), .IN4(n808), .QN(n777) );
  AOI221X1 U2595 ( .IN1(n166), .IN2(\ram[201][0] ), .IN3(n151), .IN4(
        \ram[206][0] ), .IN5(n809), .QN(n808) );
  AO22X1 U2596 ( .IN1(n769), .IN2(\ram[0][0] ), .IN3(n154), .IN4(\ram[205][0] ), .Q(n809) );
  AOI221X1 U2597 ( .IN1(n190), .IN2(\ram[193][0] ), .IN3(n175), .IN4(
        \ram[198][0] ), .IN5(n810), .QN(n807) );
  AO22X1 U2598 ( .IN1(n163), .IN2(\ram[202][0] ), .IN3(n178), .IN4(
        \ram[197][0] ), .Q(n810) );
  AOI221X1 U2599 ( .IN1(n106), .IN2(\ram[221][0] ), .IN3(n187), .IN4(
        \ram[194][0] ), .IN5(n811), .QN(n806) );
  AO22X1 U2600 ( .IN1(n103), .IN2(\ram[222][0] ), .IN3(n118), .IN4(
        \ram[217][0] ), .Q(n811) );
  AOI221X1 U2601 ( .IN1(n142), .IN2(\ram[209][0] ), .IN3(n127), .IN4(
        \ram[214][0] ), .IN5(n812), .QN(n805) );
  AO22X1 U2602 ( .IN1(n115), .IN2(\ram[218][0] ), .IN3(n130), .IN4(
        \ram[213][0] ), .Q(n812) );
  NAND4X0 U2604 ( .IN1(n817), .IN2(n818), .IN3(n819), .IN4(n820), .QN(n816) );
  AOI221X1 U2605 ( .IN1(n643), .IN2(\ram[42][0] ), .IN3(n646), .IN4(
        \ram[41][0] ), .IN5(n821), .QN(n820) );
  AO22X1 U2606 ( .IN1(n634), .IN2(\ram[45][0] ), .IN3(n631), .IN4(\ram[46][0] ), .Q(n821) );
  AOI221X1 U2607 ( .IN1(n667), .IN2(\ram[34][0] ), .IN3(n670), .IN4(
        \ram[33][0] ), .IN5(n822), .QN(n819) );
  AO22X1 U2608 ( .IN1(n658), .IN2(\ram[37][0] ), .IN3(n655), .IN4(\ram[38][0] ), .Q(n822) );
  AOI221X1 U2609 ( .IN1(n595), .IN2(\ram[58][0] ), .IN3(n598), .IN4(
        \ram[57][0] ), .IN5(n823), .QN(n818) );
  AO22X1 U2610 ( .IN1(n586), .IN2(\ram[61][0] ), .IN3(n583), .IN4(\ram[62][0] ), .Q(n823) );
  AOI221X1 U2611 ( .IN1(n619), .IN2(\ram[50][0] ), .IN3(n622), .IN4(
        \ram[49][0] ), .IN5(n824), .QN(n817) );
  AO22X1 U2612 ( .IN1(n610), .IN2(\ram[53][0] ), .IN3(n607), .IN4(\ram[54][0] ), .Q(n824) );
  NAND4X0 U2613 ( .IN1(n825), .IN2(n826), .IN3(n827), .IN4(n828), .QN(n815) );
  AOI221X1 U2614 ( .IN1(n739), .IN2(\ram[10][0] ), .IN3(n742), .IN4(
        \ram[9][0] ), .IN5(n829), .QN(n828) );
  AO22X1 U2615 ( .IN1(n730), .IN2(\ram[13][0] ), .IN3(n727), .IN4(\ram[14][0] ), .Q(n829) );
  AOI221X1 U2616 ( .IN1(n763), .IN2(\ram[2][0] ), .IN3(n766), .IN4(\ram[1][0] ), .IN5(n830), .QN(n827) );
  AO22X1 U2617 ( .IN1(n754), .IN2(\ram[5][0] ), .IN3(n751), .IN4(\ram[6][0] ), 
        .Q(n830) );
  AOI221X1 U2618 ( .IN1(n691), .IN2(\ram[26][0] ), .IN3(n694), .IN4(
        \ram[25][0] ), .IN5(n831), .QN(n826) );
  AO22X1 U2619 ( .IN1(n682), .IN2(\ram[29][0] ), .IN3(n679), .IN4(\ram[30][0] ), .Q(n831) );
  AOI221X1 U2620 ( .IN1(n715), .IN2(\ram[18][0] ), .IN3(n718), .IN4(
        \ram[17][0] ), .IN5(n832), .QN(n825) );
  AO22X1 U2621 ( .IN1(n706), .IN2(\ram[21][0] ), .IN3(n703), .IN4(\ram[22][0] ), .Q(n832) );
  NAND4X0 U2622 ( .IN1(n833), .IN2(n834), .IN3(n835), .IN4(n836), .QN(n814) );
  AOI221X1 U2623 ( .IN1(n451), .IN2(\ram[106][0] ), .IN3(n454), .IN4(
        \ram[105][0] ), .IN5(n837), .QN(n836) );
  AO22X1 U2624 ( .IN1(n442), .IN2(\ram[109][0] ), .IN3(n439), .IN4(
        \ram[110][0] ), .Q(n837) );
  AOI221X1 U2625 ( .IN1(n475), .IN2(\ram[98][0] ), .IN3(n478), .IN4(
        \ram[97][0] ), .IN5(n838), .QN(n835) );
  AO22X1 U2626 ( .IN1(n466), .IN2(\ram[101][0] ), .IN3(n463), .IN4(
        \ram[102][0] ), .Q(n838) );
  AOI221X1 U2627 ( .IN1(n403), .IN2(\ram[122][0] ), .IN3(n406), .IN4(
        \ram[121][0] ), .IN5(n839), .QN(n834) );
  AO22X1 U2628 ( .IN1(n394), .IN2(\ram[125][0] ), .IN3(n391), .IN4(
        \ram[126][0] ), .Q(n839) );
  AOI221X1 U2629 ( .IN1(n427), .IN2(\ram[114][0] ), .IN3(n430), .IN4(
        \ram[113][0] ), .IN5(n840), .QN(n833) );
  AO22X1 U2630 ( .IN1(n418), .IN2(\ram[117][0] ), .IN3(n415), .IN4(
        \ram[118][0] ), .Q(n840) );
  NAND4X0 U2631 ( .IN1(n841), .IN2(n842), .IN3(n843), .IN4(n844), .QN(n813) );
  AOI221X1 U2632 ( .IN1(n547), .IN2(\ram[74][0] ), .IN3(n550), .IN4(
        \ram[73][0] ), .IN5(n845), .QN(n844) );
  AO22X1 U2633 ( .IN1(n538), .IN2(\ram[77][0] ), .IN3(n535), .IN4(\ram[78][0] ), .Q(n845) );
  AOI221X1 U2634 ( .IN1(n571), .IN2(\ram[66][0] ), .IN3(n574), .IN4(
        \ram[65][0] ), .IN5(n846), .QN(n843) );
  AO22X1 U2635 ( .IN1(n562), .IN2(\ram[69][0] ), .IN3(n559), .IN4(\ram[70][0] ), .Q(n846) );
  AOI221X1 U2636 ( .IN1(n499), .IN2(\ram[90][0] ), .IN3(n502), .IN4(
        \ram[89][0] ), .IN5(n847), .QN(n842) );
  AO22X1 U2637 ( .IN1(n490), .IN2(\ram[93][0] ), .IN3(n487), .IN4(\ram[94][0] ), .Q(n847) );
  AOI221X1 U2638 ( .IN1(n523), .IN2(\ram[82][0] ), .IN3(n526), .IN4(
        \ram[81][0] ), .IN5(n848), .QN(n841) );
  AO22X1 U2639 ( .IN1(n514), .IN2(\ram[85][0] ), .IN3(n511), .IN4(\ram[86][0] ), .Q(n848) );
  NAND4X0 U2641 ( .IN1(n853), .IN2(n854), .IN3(n855), .IN4(n856), .QN(n852) );
  AOI221X1 U2642 ( .IN1(n253), .IN2(\ram[172][0] ), .IN3(n256), .IN4(
        \ram[171][0] ), .IN5(n857), .QN(n856) );
  AO22X1 U2643 ( .IN1(n244), .IN2(\ram[175][0] ), .IN3(n241), .IN4(
        \ram[176][0] ), .Q(n857) );
  AOI221X1 U2644 ( .IN1(n277), .IN2(\ram[164][0] ), .IN3(n280), .IN4(
        \ram[163][0] ), .IN5(n858), .QN(n855) );
  AO22X1 U2645 ( .IN1(n268), .IN2(\ram[167][0] ), .IN3(n265), .IN4(
        \ram[168][0] ), .Q(n858) );
  AOI221X1 U2646 ( .IN1(n205), .IN2(\ram[188][0] ), .IN3(n208), .IN4(
        \ram[187][0] ), .IN5(n859), .QN(n854) );
  AO22X1 U2647 ( .IN1(n202), .IN2(\ram[189][0] ), .IN3(n199), .IN4(
        \ram[190][0] ), .Q(n859) );
  AOI221X1 U2648 ( .IN1(n229), .IN2(\ram[180][0] ), .IN3(n232), .IN4(
        \ram[179][0] ), .IN5(n860), .QN(n853) );
  AO22X1 U2649 ( .IN1(n220), .IN2(\ram[183][0] ), .IN3(n217), .IN4(
        \ram[184][0] ), .Q(n860) );
  NAND4X0 U2650 ( .IN1(n861), .IN2(n862), .IN3(n863), .IN4(n864), .QN(n851) );
  AOI221X1 U2651 ( .IN1(n349), .IN2(\ram[140][0] ), .IN3(n352), .IN4(
        \ram[139][0] ), .IN5(n865), .QN(n864) );
  AO22X1 U2652 ( .IN1(n340), .IN2(\ram[143][0] ), .IN3(n337), .IN4(
        \ram[144][0] ), .Q(n865) );
  AOI221X1 U2653 ( .IN1(n373), .IN2(\ram[132][0] ), .IN3(n376), .IN4(
        \ram[131][0] ), .IN5(n866), .QN(n863) );
  AO22X1 U2654 ( .IN1(n364), .IN2(\ram[135][0] ), .IN3(n361), .IN4(
        \ram[136][0] ), .Q(n866) );
  AOI221X1 U2655 ( .IN1(n301), .IN2(\ram[156][0] ), .IN3(n304), .IN4(
        \ram[155][0] ), .IN5(n867), .QN(n862) );
  AO22X1 U2656 ( .IN1(n292), .IN2(\ram[159][0] ), .IN3(n289), .IN4(
        \ram[160][0] ), .Q(n867) );
  AOI221X1 U2657 ( .IN1(n325), .IN2(\ram[148][0] ), .IN3(n328), .IN4(
        \ram[147][0] ), .IN5(n868), .QN(n861) );
  AO22X1 U2658 ( .IN1(n316), .IN2(\ram[151][0] ), .IN3(n313), .IN4(
        \ram[152][0] ), .Q(n868) );
  NAND4X0 U2659 ( .IN1(n869), .IN2(n870), .IN3(n871), .IN4(n872), .QN(n850) );
  AOI221X1 U2660 ( .IN1(n61), .IN2(\ram[236][0] ), .IN3(n64), .IN4(
        \ram[235][0] ), .IN5(n873), .QN(n872) );
  AO22X1 U2661 ( .IN1(n58), .IN2(\ram[237][0] ), .IN3(n55), .IN4(\ram[238][0] ), .Q(n873) );
  AOI221X1 U2662 ( .IN1(n85), .IN2(\ram[228][0] ), .IN3(n88), .IN4(
        \ram[227][0] ), .IN5(n874), .QN(n871) );
  AO22X1 U2663 ( .IN1(n76), .IN2(\ram[231][0] ), .IN3(n73), .IN4(\ram[232][0] ), .Q(n874) );
  AOI221X1 U2664 ( .IN1(n19), .IN2(\ram[250][0] ), .IN3(n22), .IN4(
        \ram[249][0] ), .IN5(n875), .QN(n870) );
  AO22X1 U2665 ( .IN1(n10), .IN2(\ram[253][0] ), .IN3(n7), .IN4(\ram[254][0] ), 
        .Q(n875) );
  AOI221X1 U2666 ( .IN1(n37), .IN2(\ram[244][0] ), .IN3(n40), .IN4(
        \ram[243][0] ), .IN5(n876), .QN(n869) );
  AO22X1 U2667 ( .IN1(n28), .IN2(\ram[247][0] ), .IN3(n25), .IN4(\ram[248][0] ), .Q(n876) );
  NAND4X0 U2668 ( .IN1(n877), .IN2(n878), .IN3(n879), .IN4(n880), .QN(n849) );
  AOI221X1 U2669 ( .IN1(n157), .IN2(\ram[204][0] ), .IN3(n160), .IN4(
        \ram[203][0] ), .IN5(n881), .QN(n880) );
  AO22X1 U2670 ( .IN1(n148), .IN2(\ram[207][0] ), .IN3(n145), .IN4(
        \ram[208][0] ), .Q(n881) );
  AOI221X1 U2671 ( .IN1(n181), .IN2(\ram[196][0] ), .IN3(n184), .IN4(
        \ram[195][0] ), .IN5(n882), .QN(n879) );
  AO22X1 U2672 ( .IN1(n172), .IN2(\ram[199][0] ), .IN3(n169), .IN4(
        \ram[200][0] ), .Q(n882) );
  AOI221X1 U2673 ( .IN1(n109), .IN2(\ram[220][0] ), .IN3(n112), .IN4(
        \ram[219][0] ), .IN5(n883), .QN(n878) );
  AO22X1 U2674 ( .IN1(n100), .IN2(\ram[223][0] ), .IN3(n97), .IN4(
        \ram[224][0] ), .Q(n883) );
  AOI221X1 U2675 ( .IN1(n133), .IN2(\ram[212][0] ), .IN3(n136), .IN4(
        \ram[211][0] ), .IN5(n884), .QN(n877) );
  AO22X1 U2676 ( .IN1(n124), .IN2(\ram[215][0] ), .IN3(n121), .IN4(
        \ram[216][0] ), .Q(n884) );
  NAND4X0 U2678 ( .IN1(n889), .IN2(n890), .IN3(n891), .IN4(n892), .QN(n888) );
  AOI221X1 U2679 ( .IN1(n637), .IN2(\ram[44][0] ), .IN3(n640), .IN4(
        \ram[43][0] ), .IN5(n893), .QN(n892) );
  AO22X1 U2680 ( .IN1(n628), .IN2(\ram[47][0] ), .IN3(n625), .IN4(\ram[48][0] ), .Q(n893) );
  AOI221X1 U2681 ( .IN1(n661), .IN2(\ram[36][0] ), .IN3(n664), .IN4(
        \ram[35][0] ), .IN5(n894), .QN(n891) );
  AO22X1 U2682 ( .IN1(n652), .IN2(\ram[39][0] ), .IN3(n649), .IN4(\ram[40][0] ), .Q(n894) );
  AOI221X1 U2683 ( .IN1(n589), .IN2(\ram[60][0] ), .IN3(n592), .IN4(
        \ram[59][0] ), .IN5(n895), .QN(n890) );
  AO22X1 U2684 ( .IN1(n580), .IN2(\ram[63][0] ), .IN3(n577), .IN4(\ram[64][0] ), .Q(n895) );
  AOI221X1 U2685 ( .IN1(n613), .IN2(\ram[52][0] ), .IN3(n616), .IN4(
        \ram[51][0] ), .IN5(n896), .QN(n889) );
  AO22X1 U2686 ( .IN1(n604), .IN2(\ram[55][0] ), .IN3(n601), .IN4(\ram[56][0] ), .Q(n896) );
  NAND4X0 U2687 ( .IN1(n897), .IN2(n898), .IN3(n899), .IN4(n900), .QN(n887) );
  AOI221X1 U2688 ( .IN1(n733), .IN2(\ram[12][0] ), .IN3(n736), .IN4(
        \ram[11][0] ), .IN5(n901), .QN(n900) );
  AO22X1 U2689 ( .IN1(n724), .IN2(\ram[15][0] ), .IN3(n721), .IN4(\ram[16][0] ), .Q(n901) );
  AOI221X1 U2690 ( .IN1(n757), .IN2(\ram[4][0] ), .IN3(n760), .IN4(\ram[3][0] ), .IN5(n902), .QN(n899) );
  AO22X1 U2691 ( .IN1(n748), .IN2(\ram[7][0] ), .IN3(n745), .IN4(\ram[8][0] ), 
        .Q(n902) );
  AOI221X1 U2692 ( .IN1(n685), .IN2(\ram[28][0] ), .IN3(n688), .IN4(
        \ram[27][0] ), .IN5(n903), .QN(n898) );
  AO22X1 U2693 ( .IN1(n676), .IN2(\ram[31][0] ), .IN3(n673), .IN4(\ram[32][0] ), .Q(n903) );
  AOI221X1 U2694 ( .IN1(n709), .IN2(\ram[20][0] ), .IN3(n712), .IN4(
        \ram[19][0] ), .IN5(n904), .QN(n897) );
  AO22X1 U2695 ( .IN1(n700), .IN2(\ram[23][0] ), .IN3(n697), .IN4(\ram[24][0] ), .Q(n904) );
  NAND4X0 U2696 ( .IN1(n905), .IN2(n906), .IN3(n907), .IN4(n908), .QN(n886) );
  AOI221X1 U2697 ( .IN1(n445), .IN2(\ram[108][0] ), .IN3(n448), .IN4(
        \ram[107][0] ), .IN5(n909), .QN(n908) );
  AO22X1 U2698 ( .IN1(n436), .IN2(\ram[111][0] ), .IN3(n433), .IN4(
        \ram[112][0] ), .Q(n909) );
  AOI221X1 U2699 ( .IN1(n469), .IN2(\ram[100][0] ), .IN3(n472), .IN4(
        \ram[99][0] ), .IN5(n910), .QN(n907) );
  AO22X1 U2700 ( .IN1(n460), .IN2(\ram[103][0] ), .IN3(n457), .IN4(
        \ram[104][0] ), .Q(n910) );
  AOI221X1 U2701 ( .IN1(n397), .IN2(\ram[124][0] ), .IN3(n400), .IN4(
        \ram[123][0] ), .IN5(n911), .QN(n906) );
  AO22X1 U2702 ( .IN1(n388), .IN2(\ram[127][0] ), .IN3(n385), .IN4(
        \ram[128][0] ), .Q(n911) );
  AOI221X1 U2703 ( .IN1(n421), .IN2(\ram[116][0] ), .IN3(n424), .IN4(
        \ram[115][0] ), .IN5(n912), .QN(n905) );
  AO22X1 U2704 ( .IN1(n412), .IN2(\ram[119][0] ), .IN3(n409), .IN4(
        \ram[120][0] ), .Q(n912) );
  NAND4X0 U2705 ( .IN1(n913), .IN2(n914), .IN3(n915), .IN4(n916), .QN(n885) );
  AOI221X1 U2706 ( .IN1(n541), .IN2(\ram[76][0] ), .IN3(n544), .IN4(
        \ram[75][0] ), .IN5(n917), .QN(n916) );
  AO22X1 U2707 ( .IN1(n532), .IN2(\ram[79][0] ), .IN3(n529), .IN4(\ram[80][0] ), .Q(n917) );
  AOI221X1 U2708 ( .IN1(n565), .IN2(\ram[68][0] ), .IN3(n568), .IN4(
        \ram[67][0] ), .IN5(n918), .QN(n915) );
  AO22X1 U2709 ( .IN1(n556), .IN2(\ram[71][0] ), .IN3(n553), .IN4(\ram[72][0] ), .Q(n918) );
  AOI221X1 U2710 ( .IN1(n493), .IN2(\ram[92][0] ), .IN3(n496), .IN4(
        \ram[91][0] ), .IN5(n919), .QN(n914) );
  AO22X1 U2711 ( .IN1(n484), .IN2(\ram[95][0] ), .IN3(n481), .IN4(\ram[96][0] ), .Q(n919) );
  AOI221X1 U2712 ( .IN1(n517), .IN2(\ram[84][0] ), .IN3(n520), .IN4(
        \ram[83][0] ), .IN5(n920), .QN(n913) );
  AO22X1 U2713 ( .IN1(n508), .IN2(\ram[87][0] ), .IN3(n505), .IN4(\ram[88][0] ), .Q(n920) );
  AO22X1 U2714 ( .IN1(n771), .IN2(dataout[1]), .IN3(n4174), .IN4(n921), .Q(
        n2021) );
  NAND4X0 U2715 ( .IN1(n922), .IN2(n923), .IN3(n924), .IN4(n925), .QN(n921) );
  NAND4X0 U2717 ( .IN1(n930), .IN2(n931), .IN3(n932), .IN4(n933), .QN(n929) );
  AOI221X1 U2718 ( .IN1(n259), .IN2(\ram[170][1] ), .IN3(n262), .IN4(
        \ram[169][1] ), .IN5(n934), .QN(n933) );
  AO22X1 U2719 ( .IN1(n250), .IN2(\ram[173][1] ), .IN3(n247), .IN4(
        \ram[174][1] ), .Q(n934) );
  AOI221X1 U2720 ( .IN1(n283), .IN2(\ram[162][1] ), .IN3(n286), .IN4(
        \ram[161][1] ), .IN5(n935), .QN(n932) );
  AO22X1 U2721 ( .IN1(n274), .IN2(\ram[165][1] ), .IN3(n271), .IN4(
        \ram[166][1] ), .Q(n935) );
  AOI221X1 U2722 ( .IN1(n211), .IN2(\ram[186][1] ), .IN3(n214), .IN4(
        \ram[185][1] ), .IN5(n936), .QN(n931) );
  AO22X1 U2723 ( .IN1(n196), .IN2(\ram[191][1] ), .IN3(n193), .IN4(
        \ram[192][1] ), .Q(n936) );
  AOI221X1 U2724 ( .IN1(n235), .IN2(\ram[178][1] ), .IN3(n238), .IN4(
        \ram[177][1] ), .IN5(n937), .QN(n930) );
  AO22X1 U2725 ( .IN1(n226), .IN2(\ram[181][1] ), .IN3(n223), .IN4(
        \ram[182][1] ), .Q(n937) );
  NAND4X0 U2726 ( .IN1(n938), .IN2(n939), .IN3(n940), .IN4(n941), .QN(n928) );
  AOI221X1 U2727 ( .IN1(n355), .IN2(\ram[138][1] ), .IN3(n358), .IN4(
        \ram[137][1] ), .IN5(n942), .QN(n941) );
  AO22X1 U2728 ( .IN1(n346), .IN2(\ram[141][1] ), .IN3(n343), .IN4(
        \ram[142][1] ), .Q(n942) );
  AOI221X1 U2729 ( .IN1(n379), .IN2(\ram[130][1] ), .IN3(n382), .IN4(
        \ram[129][1] ), .IN5(n943), .QN(n940) );
  AO22X1 U2730 ( .IN1(n370), .IN2(\ram[133][1] ), .IN3(n367), .IN4(
        \ram[134][1] ), .Q(n943) );
  AOI221X1 U2731 ( .IN1(n307), .IN2(\ram[154][1] ), .IN3(n310), .IN4(
        \ram[153][1] ), .IN5(n944), .QN(n939) );
  AO22X1 U2732 ( .IN1(n298), .IN2(\ram[157][1] ), .IN3(n295), .IN4(
        \ram[158][1] ), .Q(n944) );
  AOI221X1 U2733 ( .IN1(n331), .IN2(\ram[146][1] ), .IN3(n334), .IN4(
        \ram[145][1] ), .IN5(n945), .QN(n938) );
  AO22X1 U2734 ( .IN1(n322), .IN2(\ram[149][1] ), .IN3(n319), .IN4(
        \ram[150][1] ), .Q(n945) );
  NAND4X0 U2735 ( .IN1(n946), .IN2(n947), .IN3(n948), .IN4(n949), .QN(n927) );
  AOI221X1 U2736 ( .IN1(n70), .IN2(\ram[233][1] ), .IN3(n49), .IN4(
        \ram[240][1] ), .IN5(n950), .QN(n949) );
  AO22X1 U2737 ( .IN1(n139), .IN2(\ram[210][1] ), .IN3(n52), .IN4(
        \ram[239][1] ), .Q(n950) );
  AOI221X1 U2738 ( .IN1(n94), .IN2(\ram[225][1] ), .IN3(n79), .IN4(
        \ram[230][1] ), .IN5(n951), .QN(n948) );
  AO22X1 U2739 ( .IN1(n67), .IN2(\ram[234][1] ), .IN3(n82), .IN4(\ram[229][1] ), .Q(n951) );
  AOI221X1 U2740 ( .IN1(n13), .IN2(\ram[252][1] ), .IN3(n16), .IN4(
        \ram[251][1] ), .IN5(n952), .QN(n947) );
  AO22X1 U2741 ( .IN1(n91), .IN2(\ram[226][1] ), .IN3(n3), .IN4(\ram[255][1] ), 
        .Q(n952) );
  AOI221X1 U2742 ( .IN1(n43), .IN2(\ram[242][1] ), .IN3(n46), .IN4(
        \ram[241][1] ), .IN5(n953), .QN(n946) );
  AO22X1 U2743 ( .IN1(n34), .IN2(\ram[245][1] ), .IN3(n31), .IN4(\ram[246][1] ), .Q(n953) );
  NAND4X0 U2744 ( .IN1(n954), .IN2(n955), .IN3(n956), .IN4(n957), .QN(n926) );
  AOI221X1 U2745 ( .IN1(n166), .IN2(\ram[201][1] ), .IN3(n151), .IN4(
        \ram[206][1] ), .IN5(n958), .QN(n957) );
  AO22X1 U2746 ( .IN1(n769), .IN2(\ram[0][1] ), .IN3(n154), .IN4(\ram[205][1] ), .Q(n958) );
  AOI221X1 U2747 ( .IN1(n190), .IN2(\ram[193][1] ), .IN3(n175), .IN4(
        \ram[198][1] ), .IN5(n959), .QN(n956) );
  AO22X1 U2748 ( .IN1(n163), .IN2(\ram[202][1] ), .IN3(n178), .IN4(
        \ram[197][1] ), .Q(n959) );
  AOI221X1 U2749 ( .IN1(n106), .IN2(\ram[221][1] ), .IN3(n187), .IN4(
        \ram[194][1] ), .IN5(n960), .QN(n955) );
  AO22X1 U2750 ( .IN1(n103), .IN2(\ram[222][1] ), .IN3(n118), .IN4(
        \ram[217][1] ), .Q(n960) );
  AOI221X1 U2751 ( .IN1(n142), .IN2(\ram[209][1] ), .IN3(n127), .IN4(
        \ram[214][1] ), .IN5(n961), .QN(n954) );
  AO22X1 U2752 ( .IN1(n115), .IN2(\ram[218][1] ), .IN3(n130), .IN4(
        \ram[213][1] ), .Q(n961) );
  NAND4X0 U2754 ( .IN1(n966), .IN2(n967), .IN3(n968), .IN4(n969), .QN(n965) );
  AOI221X1 U2755 ( .IN1(n643), .IN2(\ram[42][1] ), .IN3(n646), .IN4(
        \ram[41][1] ), .IN5(n970), .QN(n969) );
  AO22X1 U2756 ( .IN1(n634), .IN2(\ram[45][1] ), .IN3(n631), .IN4(\ram[46][1] ), .Q(n970) );
  AOI221X1 U2757 ( .IN1(n667), .IN2(\ram[34][1] ), .IN3(n670), .IN4(
        \ram[33][1] ), .IN5(n971), .QN(n968) );
  AO22X1 U2758 ( .IN1(n658), .IN2(\ram[37][1] ), .IN3(n655), .IN4(\ram[38][1] ), .Q(n971) );
  AOI221X1 U2759 ( .IN1(n595), .IN2(\ram[58][1] ), .IN3(n598), .IN4(
        \ram[57][1] ), .IN5(n972), .QN(n967) );
  AO22X1 U2760 ( .IN1(n586), .IN2(\ram[61][1] ), .IN3(n583), .IN4(\ram[62][1] ), .Q(n972) );
  AOI221X1 U2761 ( .IN1(n619), .IN2(\ram[50][1] ), .IN3(n622), .IN4(
        \ram[49][1] ), .IN5(n973), .QN(n966) );
  AO22X1 U2762 ( .IN1(n610), .IN2(\ram[53][1] ), .IN3(n607), .IN4(\ram[54][1] ), .Q(n973) );
  NAND4X0 U2763 ( .IN1(n974), .IN2(n975), .IN3(n976), .IN4(n977), .QN(n964) );
  AOI221X1 U2764 ( .IN1(n739), .IN2(\ram[10][1] ), .IN3(n742), .IN4(
        \ram[9][1] ), .IN5(n978), .QN(n977) );
  AO22X1 U2765 ( .IN1(n730), .IN2(\ram[13][1] ), .IN3(n727), .IN4(\ram[14][1] ), .Q(n978) );
  AOI221X1 U2766 ( .IN1(n763), .IN2(\ram[2][1] ), .IN3(n766), .IN4(\ram[1][1] ), .IN5(n979), .QN(n976) );
  AO22X1 U2767 ( .IN1(n754), .IN2(\ram[5][1] ), .IN3(n751), .IN4(\ram[6][1] ), 
        .Q(n979) );
  AOI221X1 U2768 ( .IN1(n691), .IN2(\ram[26][1] ), .IN3(n694), .IN4(
        \ram[25][1] ), .IN5(n980), .QN(n975) );
  AO22X1 U2769 ( .IN1(n682), .IN2(\ram[29][1] ), .IN3(n679), .IN4(\ram[30][1] ), .Q(n980) );
  AOI221X1 U2770 ( .IN1(n715), .IN2(\ram[18][1] ), .IN3(n718), .IN4(
        \ram[17][1] ), .IN5(n981), .QN(n974) );
  AO22X1 U2771 ( .IN1(n706), .IN2(\ram[21][1] ), .IN3(n703), .IN4(\ram[22][1] ), .Q(n981) );
  NAND4X0 U2772 ( .IN1(n982), .IN2(n983), .IN3(n984), .IN4(n985), .QN(n963) );
  AOI221X1 U2773 ( .IN1(n451), .IN2(\ram[106][1] ), .IN3(n454), .IN4(
        \ram[105][1] ), .IN5(n986), .QN(n985) );
  AO22X1 U2774 ( .IN1(n442), .IN2(\ram[109][1] ), .IN3(n439), .IN4(
        \ram[110][1] ), .Q(n986) );
  AOI221X1 U2775 ( .IN1(n475), .IN2(\ram[98][1] ), .IN3(n478), .IN4(
        \ram[97][1] ), .IN5(n987), .QN(n984) );
  AO22X1 U2776 ( .IN1(n466), .IN2(\ram[101][1] ), .IN3(n463), .IN4(
        \ram[102][1] ), .Q(n987) );
  AOI221X1 U2777 ( .IN1(n403), .IN2(\ram[122][1] ), .IN3(n406), .IN4(
        \ram[121][1] ), .IN5(n988), .QN(n983) );
  AO22X1 U2778 ( .IN1(n394), .IN2(\ram[125][1] ), .IN3(n391), .IN4(
        \ram[126][1] ), .Q(n988) );
  AOI221X1 U2779 ( .IN1(n427), .IN2(\ram[114][1] ), .IN3(n430), .IN4(
        \ram[113][1] ), .IN5(n989), .QN(n982) );
  AO22X1 U2780 ( .IN1(n418), .IN2(\ram[117][1] ), .IN3(n415), .IN4(
        \ram[118][1] ), .Q(n989) );
  NAND4X0 U2781 ( .IN1(n990), .IN2(n991), .IN3(n992), .IN4(n993), .QN(n962) );
  AOI221X1 U2782 ( .IN1(n547), .IN2(\ram[74][1] ), .IN3(n550), .IN4(
        \ram[73][1] ), .IN5(n994), .QN(n993) );
  AO22X1 U2783 ( .IN1(n538), .IN2(\ram[77][1] ), .IN3(n535), .IN4(\ram[78][1] ), .Q(n994) );
  AOI221X1 U2784 ( .IN1(n571), .IN2(\ram[66][1] ), .IN3(n574), .IN4(
        \ram[65][1] ), .IN5(n995), .QN(n992) );
  AO22X1 U2785 ( .IN1(n562), .IN2(\ram[69][1] ), .IN3(n559), .IN4(\ram[70][1] ), .Q(n995) );
  AOI221X1 U2786 ( .IN1(n499), .IN2(\ram[90][1] ), .IN3(n502), .IN4(
        \ram[89][1] ), .IN5(n996), .QN(n991) );
  AO22X1 U2787 ( .IN1(n490), .IN2(\ram[93][1] ), .IN3(n487), .IN4(\ram[94][1] ), .Q(n996) );
  AOI221X1 U2788 ( .IN1(n523), .IN2(\ram[82][1] ), .IN3(n526), .IN4(
        \ram[81][1] ), .IN5(n997), .QN(n990) );
  AO22X1 U2789 ( .IN1(n514), .IN2(\ram[85][1] ), .IN3(n511), .IN4(\ram[86][1] ), .Q(n997) );
  NAND4X0 U2791 ( .IN1(n1002), .IN2(n1003), .IN3(n1004), .IN4(n1005), .QN(
        n1001) );
  AOI221X1 U2792 ( .IN1(n253), .IN2(\ram[172][1] ), .IN3(n256), .IN4(
        \ram[171][1] ), .IN5(n1006), .QN(n1005) );
  AO22X1 U2793 ( .IN1(n244), .IN2(\ram[175][1] ), .IN3(n241), .IN4(
        \ram[176][1] ), .Q(n1006) );
  AOI221X1 U2794 ( .IN1(n277), .IN2(\ram[164][1] ), .IN3(n280), .IN4(
        \ram[163][1] ), .IN5(n1007), .QN(n1004) );
  AO22X1 U2795 ( .IN1(n268), .IN2(\ram[167][1] ), .IN3(n265), .IN4(
        \ram[168][1] ), .Q(n1007) );
  AOI221X1 U2796 ( .IN1(n205), .IN2(\ram[188][1] ), .IN3(n208), .IN4(
        \ram[187][1] ), .IN5(n1008), .QN(n1003) );
  AO22X1 U2797 ( .IN1(n202), .IN2(\ram[189][1] ), .IN3(n199), .IN4(
        \ram[190][1] ), .Q(n1008) );
  AOI221X1 U2798 ( .IN1(n229), .IN2(\ram[180][1] ), .IN3(n232), .IN4(
        \ram[179][1] ), .IN5(n1009), .QN(n1002) );
  AO22X1 U2799 ( .IN1(n220), .IN2(\ram[183][1] ), .IN3(n217), .IN4(
        \ram[184][1] ), .Q(n1009) );
  NAND4X0 U2800 ( .IN1(n1010), .IN2(n1011), .IN3(n1012), .IN4(n1013), .QN(
        n1000) );
  AOI221X1 U2801 ( .IN1(n349), .IN2(\ram[140][1] ), .IN3(n352), .IN4(
        \ram[139][1] ), .IN5(n1014), .QN(n1013) );
  AO22X1 U2802 ( .IN1(n340), .IN2(\ram[143][1] ), .IN3(n337), .IN4(
        \ram[144][1] ), .Q(n1014) );
  AOI221X1 U2803 ( .IN1(n373), .IN2(\ram[132][1] ), .IN3(n376), .IN4(
        \ram[131][1] ), .IN5(n1015), .QN(n1012) );
  AO22X1 U2804 ( .IN1(n364), .IN2(\ram[135][1] ), .IN3(n361), .IN4(
        \ram[136][1] ), .Q(n1015) );
  AOI221X1 U2805 ( .IN1(n301), .IN2(\ram[156][1] ), .IN3(n304), .IN4(
        \ram[155][1] ), .IN5(n1016), .QN(n1011) );
  AO22X1 U2806 ( .IN1(n292), .IN2(\ram[159][1] ), .IN3(n289), .IN4(
        \ram[160][1] ), .Q(n1016) );
  AOI221X1 U2807 ( .IN1(n325), .IN2(\ram[148][1] ), .IN3(n328), .IN4(
        \ram[147][1] ), .IN5(n1017), .QN(n1010) );
  AO22X1 U2808 ( .IN1(n316), .IN2(\ram[151][1] ), .IN3(n313), .IN4(
        \ram[152][1] ), .Q(n1017) );
  NAND4X0 U2809 ( .IN1(n1018), .IN2(n1019), .IN3(n1020), .IN4(n1021), .QN(n999) );
  AOI221X1 U2810 ( .IN1(n61), .IN2(\ram[236][1] ), .IN3(n64), .IN4(
        \ram[235][1] ), .IN5(n1022), .QN(n1021) );
  AO22X1 U2811 ( .IN1(n58), .IN2(\ram[237][1] ), .IN3(n55), .IN4(\ram[238][1] ), .Q(n1022) );
  AOI221X1 U2812 ( .IN1(n85), .IN2(\ram[228][1] ), .IN3(n88), .IN4(
        \ram[227][1] ), .IN5(n1023), .QN(n1020) );
  AO22X1 U2813 ( .IN1(n76), .IN2(\ram[231][1] ), .IN3(n73), .IN4(\ram[232][1] ), .Q(n1023) );
  AOI221X1 U2814 ( .IN1(n19), .IN2(\ram[250][1] ), .IN3(n22), .IN4(
        \ram[249][1] ), .IN5(n1024), .QN(n1019) );
  AO22X1 U2815 ( .IN1(n10), .IN2(\ram[253][1] ), .IN3(n7), .IN4(\ram[254][1] ), 
        .Q(n1024) );
  AOI221X1 U2816 ( .IN1(n37), .IN2(\ram[244][1] ), .IN3(n40), .IN4(
        \ram[243][1] ), .IN5(n1025), .QN(n1018) );
  AO22X1 U2817 ( .IN1(n28), .IN2(\ram[247][1] ), .IN3(n25), .IN4(\ram[248][1] ), .Q(n1025) );
  NAND4X0 U2818 ( .IN1(n1026), .IN2(n1027), .IN3(n1028), .IN4(n1029), .QN(n998) );
  AOI221X1 U2819 ( .IN1(n157), .IN2(\ram[204][1] ), .IN3(n160), .IN4(
        \ram[203][1] ), .IN5(n1030), .QN(n1029) );
  AO22X1 U2820 ( .IN1(n148), .IN2(\ram[207][1] ), .IN3(n145), .IN4(
        \ram[208][1] ), .Q(n1030) );
  AOI221X1 U2821 ( .IN1(n181), .IN2(\ram[196][1] ), .IN3(n184), .IN4(
        \ram[195][1] ), .IN5(n1031), .QN(n1028) );
  AO22X1 U2822 ( .IN1(n172), .IN2(\ram[199][1] ), .IN3(n169), .IN4(
        \ram[200][1] ), .Q(n1031) );
  AOI221X1 U2823 ( .IN1(n109), .IN2(\ram[220][1] ), .IN3(n112), .IN4(
        \ram[219][1] ), .IN5(n1032), .QN(n1027) );
  AO22X1 U2824 ( .IN1(n100), .IN2(\ram[223][1] ), .IN3(n97), .IN4(
        \ram[224][1] ), .Q(n1032) );
  AOI221X1 U2825 ( .IN1(n133), .IN2(\ram[212][1] ), .IN3(n136), .IN4(
        \ram[211][1] ), .IN5(n1033), .QN(n1026) );
  AO22X1 U2826 ( .IN1(n124), .IN2(\ram[215][1] ), .IN3(n121), .IN4(
        \ram[216][1] ), .Q(n1033) );
  NAND4X0 U2828 ( .IN1(n1038), .IN2(n1039), .IN3(n1040), .IN4(n1041), .QN(
        n1037) );
  AOI221X1 U2829 ( .IN1(n637), .IN2(\ram[44][1] ), .IN3(n640), .IN4(
        \ram[43][1] ), .IN5(n1042), .QN(n1041) );
  AO22X1 U2830 ( .IN1(n628), .IN2(\ram[47][1] ), .IN3(n625), .IN4(\ram[48][1] ), .Q(n1042) );
  AOI221X1 U2831 ( .IN1(n661), .IN2(\ram[36][1] ), .IN3(n664), .IN4(
        \ram[35][1] ), .IN5(n1043), .QN(n1040) );
  AO22X1 U2832 ( .IN1(n652), .IN2(\ram[39][1] ), .IN3(n649), .IN4(\ram[40][1] ), .Q(n1043) );
  AOI221X1 U2833 ( .IN1(n589), .IN2(\ram[60][1] ), .IN3(n592), .IN4(
        \ram[59][1] ), .IN5(n1044), .QN(n1039) );
  AO22X1 U2834 ( .IN1(n580), .IN2(\ram[63][1] ), .IN3(n577), .IN4(\ram[64][1] ), .Q(n1044) );
  AOI221X1 U2835 ( .IN1(n613), .IN2(\ram[52][1] ), .IN3(n616), .IN4(
        \ram[51][1] ), .IN5(n1045), .QN(n1038) );
  AO22X1 U2836 ( .IN1(n604), .IN2(\ram[55][1] ), .IN3(n601), .IN4(\ram[56][1] ), .Q(n1045) );
  NAND4X0 U2837 ( .IN1(n1046), .IN2(n1047), .IN3(n1048), .IN4(n1049), .QN(
        n1036) );
  AOI221X1 U2838 ( .IN1(n733), .IN2(\ram[12][1] ), .IN3(n736), .IN4(
        \ram[11][1] ), .IN5(n1050), .QN(n1049) );
  AO22X1 U2839 ( .IN1(n724), .IN2(\ram[15][1] ), .IN3(n721), .IN4(\ram[16][1] ), .Q(n1050) );
  AOI221X1 U2840 ( .IN1(n757), .IN2(\ram[4][1] ), .IN3(n760), .IN4(\ram[3][1] ), .IN5(n1051), .QN(n1048) );
  AO22X1 U2841 ( .IN1(n748), .IN2(\ram[7][1] ), .IN3(n745), .IN4(\ram[8][1] ), 
        .Q(n1051) );
  AOI221X1 U2842 ( .IN1(n685), .IN2(\ram[28][1] ), .IN3(n688), .IN4(
        \ram[27][1] ), .IN5(n1052), .QN(n1047) );
  AO22X1 U2843 ( .IN1(n676), .IN2(\ram[31][1] ), .IN3(n673), .IN4(\ram[32][1] ), .Q(n1052) );
  AOI221X1 U2844 ( .IN1(n709), .IN2(\ram[20][1] ), .IN3(n712), .IN4(
        \ram[19][1] ), .IN5(n1053), .QN(n1046) );
  AO22X1 U2845 ( .IN1(n700), .IN2(\ram[23][1] ), .IN3(n697), .IN4(\ram[24][1] ), .Q(n1053) );
  NAND4X0 U2846 ( .IN1(n1054), .IN2(n1055), .IN3(n1056), .IN4(n1057), .QN(
        n1035) );
  AOI221X1 U2847 ( .IN1(n445), .IN2(\ram[108][1] ), .IN3(n448), .IN4(
        \ram[107][1] ), .IN5(n1058), .QN(n1057) );
  AO22X1 U2848 ( .IN1(n436), .IN2(\ram[111][1] ), .IN3(n433), .IN4(
        \ram[112][1] ), .Q(n1058) );
  AOI221X1 U2849 ( .IN1(n469), .IN2(\ram[100][1] ), .IN3(n472), .IN4(
        \ram[99][1] ), .IN5(n1059), .QN(n1056) );
  AO22X1 U2850 ( .IN1(n460), .IN2(\ram[103][1] ), .IN3(n457), .IN4(
        \ram[104][1] ), .Q(n1059) );
  AOI221X1 U2851 ( .IN1(n397), .IN2(\ram[124][1] ), .IN3(n400), .IN4(
        \ram[123][1] ), .IN5(n1060), .QN(n1055) );
  AO22X1 U2852 ( .IN1(n388), .IN2(\ram[127][1] ), .IN3(n385), .IN4(
        \ram[128][1] ), .Q(n1060) );
  AOI221X1 U2853 ( .IN1(n421), .IN2(\ram[116][1] ), .IN3(n424), .IN4(
        \ram[115][1] ), .IN5(n1061), .QN(n1054) );
  AO22X1 U2854 ( .IN1(n412), .IN2(\ram[119][1] ), .IN3(n409), .IN4(
        \ram[120][1] ), .Q(n1061) );
  NAND4X0 U2855 ( .IN1(n1062), .IN2(n1063), .IN3(n1064), .IN4(n1065), .QN(
        n1034) );
  AOI221X1 U2856 ( .IN1(n541), .IN2(\ram[76][1] ), .IN3(n544), .IN4(
        \ram[75][1] ), .IN5(n1066), .QN(n1065) );
  AO22X1 U2857 ( .IN1(n532), .IN2(\ram[79][1] ), .IN3(n529), .IN4(\ram[80][1] ), .Q(n1066) );
  AOI221X1 U2858 ( .IN1(n565), .IN2(\ram[68][1] ), .IN3(n568), .IN4(
        \ram[67][1] ), .IN5(n1067), .QN(n1064) );
  AO22X1 U2859 ( .IN1(n556), .IN2(\ram[71][1] ), .IN3(n553), .IN4(\ram[72][1] ), .Q(n1067) );
  AOI221X1 U2860 ( .IN1(n493), .IN2(\ram[92][1] ), .IN3(n496), .IN4(
        \ram[91][1] ), .IN5(n1068), .QN(n1063) );
  AO22X1 U2861 ( .IN1(n484), .IN2(\ram[95][1] ), .IN3(n481), .IN4(\ram[96][1] ), .Q(n1068) );
  AOI221X1 U2862 ( .IN1(n517), .IN2(\ram[84][1] ), .IN3(n520), .IN4(
        \ram[83][1] ), .IN5(n1069), .QN(n1062) );
  AO22X1 U2863 ( .IN1(n508), .IN2(\ram[87][1] ), .IN3(n505), .IN4(\ram[88][1] ), .Q(n1069) );
  AO22X1 U2864 ( .IN1(n771), .IN2(dataout[2]), .IN3(n4174), .IN4(n1070), .Q(
        n2022) );
  NAND4X0 U2865 ( .IN1(n1071), .IN2(n1072), .IN3(n1073), .IN4(n1074), .QN(
        n1070) );
  NAND4X0 U2867 ( .IN1(n1079), .IN2(n1080), .IN3(n1081), .IN4(n1082), .QN(
        n1078) );
  AOI221X1 U2868 ( .IN1(n259), .IN2(\ram[170][2] ), .IN3(n262), .IN4(
        \ram[169][2] ), .IN5(n1083), .QN(n1082) );
  AO22X1 U2869 ( .IN1(n250), .IN2(\ram[173][2] ), .IN3(n247), .IN4(
        \ram[174][2] ), .Q(n1083) );
  AOI221X1 U2870 ( .IN1(n283), .IN2(\ram[162][2] ), .IN3(n286), .IN4(
        \ram[161][2] ), .IN5(n1084), .QN(n1081) );
  AO22X1 U2871 ( .IN1(n274), .IN2(\ram[165][2] ), .IN3(n271), .IN4(
        \ram[166][2] ), .Q(n1084) );
  AOI221X1 U2872 ( .IN1(n211), .IN2(\ram[186][2] ), .IN3(n214), .IN4(
        \ram[185][2] ), .IN5(n1085), .QN(n1080) );
  AO22X1 U2873 ( .IN1(n196), .IN2(\ram[191][2] ), .IN3(n193), .IN4(
        \ram[192][2] ), .Q(n1085) );
  AOI221X1 U2874 ( .IN1(n235), .IN2(\ram[178][2] ), .IN3(n238), .IN4(
        \ram[177][2] ), .IN5(n1086), .QN(n1079) );
  AO22X1 U2875 ( .IN1(n226), .IN2(\ram[181][2] ), .IN3(n223), .IN4(
        \ram[182][2] ), .Q(n1086) );
  NAND4X0 U2876 ( .IN1(n1087), .IN2(n1088), .IN3(n1089), .IN4(n1090), .QN(
        n1077) );
  AOI221X1 U2877 ( .IN1(n355), .IN2(\ram[138][2] ), .IN3(n358), .IN4(
        \ram[137][2] ), .IN5(n1091), .QN(n1090) );
  AO22X1 U2878 ( .IN1(n346), .IN2(\ram[141][2] ), .IN3(n343), .IN4(
        \ram[142][2] ), .Q(n1091) );
  AOI221X1 U2879 ( .IN1(n379), .IN2(\ram[130][2] ), .IN3(n382), .IN4(
        \ram[129][2] ), .IN5(n1092), .QN(n1089) );
  AO22X1 U2880 ( .IN1(n370), .IN2(\ram[133][2] ), .IN3(n367), .IN4(
        \ram[134][2] ), .Q(n1092) );
  AOI221X1 U2881 ( .IN1(n307), .IN2(\ram[154][2] ), .IN3(n310), .IN4(
        \ram[153][2] ), .IN5(n1093), .QN(n1088) );
  AO22X1 U2882 ( .IN1(n298), .IN2(\ram[157][2] ), .IN3(n295), .IN4(
        \ram[158][2] ), .Q(n1093) );
  AOI221X1 U2883 ( .IN1(n331), .IN2(\ram[146][2] ), .IN3(n334), .IN4(
        \ram[145][2] ), .IN5(n1094), .QN(n1087) );
  AO22X1 U2884 ( .IN1(n322), .IN2(\ram[149][2] ), .IN3(n319), .IN4(
        \ram[150][2] ), .Q(n1094) );
  NAND4X0 U2885 ( .IN1(n1095), .IN2(n1096), .IN3(n1097), .IN4(n1098), .QN(
        n1076) );
  AOI221X1 U2886 ( .IN1(n70), .IN2(\ram[233][2] ), .IN3(n49), .IN4(
        \ram[240][2] ), .IN5(n1099), .QN(n1098) );
  AO22X1 U2887 ( .IN1(n139), .IN2(\ram[210][2] ), .IN3(n52), .IN4(
        \ram[239][2] ), .Q(n1099) );
  AOI221X1 U2888 ( .IN1(n94), .IN2(\ram[225][2] ), .IN3(n79), .IN4(
        \ram[230][2] ), .IN5(n1100), .QN(n1097) );
  AO22X1 U2889 ( .IN1(n67), .IN2(\ram[234][2] ), .IN3(n82), .IN4(\ram[229][2] ), .Q(n1100) );
  AOI221X1 U2890 ( .IN1(n13), .IN2(\ram[252][2] ), .IN3(n16), .IN4(
        \ram[251][2] ), .IN5(n1101), .QN(n1096) );
  AO22X1 U2891 ( .IN1(n91), .IN2(\ram[226][2] ), .IN3(n3), .IN4(\ram[255][2] ), 
        .Q(n1101) );
  AOI221X1 U2892 ( .IN1(n43), .IN2(\ram[242][2] ), .IN3(n46), .IN4(
        \ram[241][2] ), .IN5(n1102), .QN(n1095) );
  AO22X1 U2893 ( .IN1(n34), .IN2(\ram[245][2] ), .IN3(n31), .IN4(\ram[246][2] ), .Q(n1102) );
  NAND4X0 U2894 ( .IN1(n1103), .IN2(n1104), .IN3(n1105), .IN4(n1106), .QN(
        n1075) );
  AOI221X1 U2895 ( .IN1(n166), .IN2(\ram[201][2] ), .IN3(n151), .IN4(
        \ram[206][2] ), .IN5(n1107), .QN(n1106) );
  AO22X1 U2896 ( .IN1(n769), .IN2(\ram[0][2] ), .IN3(n154), .IN4(\ram[205][2] ), .Q(n1107) );
  AOI221X1 U2897 ( .IN1(n190), .IN2(\ram[193][2] ), .IN3(n175), .IN4(
        \ram[198][2] ), .IN5(n1108), .QN(n1105) );
  AO22X1 U2898 ( .IN1(n163), .IN2(\ram[202][2] ), .IN3(n178), .IN4(
        \ram[197][2] ), .Q(n1108) );
  AOI221X1 U2899 ( .IN1(n106), .IN2(\ram[221][2] ), .IN3(n187), .IN4(
        \ram[194][2] ), .IN5(n1109), .QN(n1104) );
  AO22X1 U2900 ( .IN1(n103), .IN2(\ram[222][2] ), .IN3(n118), .IN4(
        \ram[217][2] ), .Q(n1109) );
  AOI221X1 U2901 ( .IN1(n142), .IN2(\ram[209][2] ), .IN3(n127), .IN4(
        \ram[214][2] ), .IN5(n1110), .QN(n1103) );
  AO22X1 U2902 ( .IN1(n115), .IN2(\ram[218][2] ), .IN3(n130), .IN4(
        \ram[213][2] ), .Q(n1110) );
  NAND4X0 U2904 ( .IN1(n1115), .IN2(n1116), .IN3(n1117), .IN4(n1118), .QN(
        n1114) );
  AOI221X1 U2905 ( .IN1(n643), .IN2(\ram[42][2] ), .IN3(n646), .IN4(
        \ram[41][2] ), .IN5(n1119), .QN(n1118) );
  AO22X1 U2906 ( .IN1(n634), .IN2(\ram[45][2] ), .IN3(n631), .IN4(\ram[46][2] ), .Q(n1119) );
  AOI221X1 U2907 ( .IN1(n667), .IN2(\ram[34][2] ), .IN3(n670), .IN4(
        \ram[33][2] ), .IN5(n1120), .QN(n1117) );
  AO22X1 U2908 ( .IN1(n658), .IN2(\ram[37][2] ), .IN3(n655), .IN4(\ram[38][2] ), .Q(n1120) );
  AOI221X1 U2909 ( .IN1(n595), .IN2(\ram[58][2] ), .IN3(n598), .IN4(
        \ram[57][2] ), .IN5(n1121), .QN(n1116) );
  AO22X1 U2910 ( .IN1(n586), .IN2(\ram[61][2] ), .IN3(n583), .IN4(\ram[62][2] ), .Q(n1121) );
  AOI221X1 U2911 ( .IN1(n619), .IN2(\ram[50][2] ), .IN3(n622), .IN4(
        \ram[49][2] ), .IN5(n1122), .QN(n1115) );
  AO22X1 U2912 ( .IN1(n610), .IN2(\ram[53][2] ), .IN3(n607), .IN4(\ram[54][2] ), .Q(n1122) );
  NAND4X0 U2913 ( .IN1(n1123), .IN2(n1124), .IN3(n1125), .IN4(n1126), .QN(
        n1113) );
  AOI221X1 U2914 ( .IN1(n739), .IN2(\ram[10][2] ), .IN3(n742), .IN4(
        \ram[9][2] ), .IN5(n1127), .QN(n1126) );
  AO22X1 U2915 ( .IN1(n730), .IN2(\ram[13][2] ), .IN3(n727), .IN4(\ram[14][2] ), .Q(n1127) );
  AOI221X1 U2916 ( .IN1(n763), .IN2(\ram[2][2] ), .IN3(n766), .IN4(\ram[1][2] ), .IN5(n1128), .QN(n1125) );
  AO22X1 U2917 ( .IN1(n754), .IN2(\ram[5][2] ), .IN3(n751), .IN4(\ram[6][2] ), 
        .Q(n1128) );
  AOI221X1 U2918 ( .IN1(n691), .IN2(\ram[26][2] ), .IN3(n694), .IN4(
        \ram[25][2] ), .IN5(n1129), .QN(n1124) );
  AO22X1 U2919 ( .IN1(n682), .IN2(\ram[29][2] ), .IN3(n679), .IN4(\ram[30][2] ), .Q(n1129) );
  AOI221X1 U2920 ( .IN1(n715), .IN2(\ram[18][2] ), .IN3(n718), .IN4(
        \ram[17][2] ), .IN5(n1130), .QN(n1123) );
  AO22X1 U2921 ( .IN1(n706), .IN2(\ram[21][2] ), .IN3(n703), .IN4(\ram[22][2] ), .Q(n1130) );
  NAND4X0 U2922 ( .IN1(n1131), .IN2(n1132), .IN3(n1133), .IN4(n1134), .QN(
        n1112) );
  AOI221X1 U2923 ( .IN1(n451), .IN2(\ram[106][2] ), .IN3(n454), .IN4(
        \ram[105][2] ), .IN5(n1135), .QN(n1134) );
  AO22X1 U2924 ( .IN1(n442), .IN2(\ram[109][2] ), .IN3(n439), .IN4(
        \ram[110][2] ), .Q(n1135) );
  AOI221X1 U2925 ( .IN1(n475), .IN2(\ram[98][2] ), .IN3(n478), .IN4(
        \ram[97][2] ), .IN5(n1136), .QN(n1133) );
  AO22X1 U2926 ( .IN1(n466), .IN2(\ram[101][2] ), .IN3(n463), .IN4(
        \ram[102][2] ), .Q(n1136) );
  AOI221X1 U2927 ( .IN1(n403), .IN2(\ram[122][2] ), .IN3(n406), .IN4(
        \ram[121][2] ), .IN5(n1137), .QN(n1132) );
  AO22X1 U2928 ( .IN1(n394), .IN2(\ram[125][2] ), .IN3(n391), .IN4(
        \ram[126][2] ), .Q(n1137) );
  AOI221X1 U2929 ( .IN1(n427), .IN2(\ram[114][2] ), .IN3(n430), .IN4(
        \ram[113][2] ), .IN5(n1138), .QN(n1131) );
  AO22X1 U2930 ( .IN1(n418), .IN2(\ram[117][2] ), .IN3(n415), .IN4(
        \ram[118][2] ), .Q(n1138) );
  NAND4X0 U2931 ( .IN1(n1139), .IN2(n1140), .IN3(n1141), .IN4(n1142), .QN(
        n1111) );
  AOI221X1 U2932 ( .IN1(n547), .IN2(\ram[74][2] ), .IN3(n550), .IN4(
        \ram[73][2] ), .IN5(n1143), .QN(n1142) );
  AO22X1 U2933 ( .IN1(n538), .IN2(\ram[77][2] ), .IN3(n535), .IN4(\ram[78][2] ), .Q(n1143) );
  AOI221X1 U2934 ( .IN1(n571), .IN2(\ram[66][2] ), .IN3(n574), .IN4(
        \ram[65][2] ), .IN5(n1144), .QN(n1141) );
  AO22X1 U2935 ( .IN1(n562), .IN2(\ram[69][2] ), .IN3(n559), .IN4(\ram[70][2] ), .Q(n1144) );
  AOI221X1 U2936 ( .IN1(n499), .IN2(\ram[90][2] ), .IN3(n502), .IN4(
        \ram[89][2] ), .IN5(n1145), .QN(n1140) );
  AO22X1 U2937 ( .IN1(n490), .IN2(\ram[93][2] ), .IN3(n487), .IN4(\ram[94][2] ), .Q(n1145) );
  AOI221X1 U2938 ( .IN1(n523), .IN2(\ram[82][2] ), .IN3(n526), .IN4(
        \ram[81][2] ), .IN5(n1146), .QN(n1139) );
  AO22X1 U2939 ( .IN1(n514), .IN2(\ram[85][2] ), .IN3(n511), .IN4(\ram[86][2] ), .Q(n1146) );
  NAND4X0 U2941 ( .IN1(n1151), .IN2(n1152), .IN3(n1153), .IN4(n1154), .QN(
        n1150) );
  AOI221X1 U2942 ( .IN1(n253), .IN2(\ram[172][2] ), .IN3(n256), .IN4(
        \ram[171][2] ), .IN5(n1155), .QN(n1154) );
  AO22X1 U2943 ( .IN1(n244), .IN2(\ram[175][2] ), .IN3(n241), .IN4(
        \ram[176][2] ), .Q(n1155) );
  AOI221X1 U2944 ( .IN1(n277), .IN2(\ram[164][2] ), .IN3(n280), .IN4(
        \ram[163][2] ), .IN5(n1156), .QN(n1153) );
  AO22X1 U2945 ( .IN1(n268), .IN2(\ram[167][2] ), .IN3(n265), .IN4(
        \ram[168][2] ), .Q(n1156) );
  AOI221X1 U2946 ( .IN1(n205), .IN2(\ram[188][2] ), .IN3(n208), .IN4(
        \ram[187][2] ), .IN5(n1157), .QN(n1152) );
  AO22X1 U2947 ( .IN1(n202), .IN2(\ram[189][2] ), .IN3(n199), .IN4(
        \ram[190][2] ), .Q(n1157) );
  AOI221X1 U2948 ( .IN1(n229), .IN2(\ram[180][2] ), .IN3(n232), .IN4(
        \ram[179][2] ), .IN5(n1158), .QN(n1151) );
  AO22X1 U2949 ( .IN1(n220), .IN2(\ram[183][2] ), .IN3(n217), .IN4(
        \ram[184][2] ), .Q(n1158) );
  NAND4X0 U2950 ( .IN1(n1159), .IN2(n1160), .IN3(n1161), .IN4(n1162), .QN(
        n1149) );
  AOI221X1 U2951 ( .IN1(n349), .IN2(\ram[140][2] ), .IN3(n352), .IN4(
        \ram[139][2] ), .IN5(n1163), .QN(n1162) );
  AO22X1 U2952 ( .IN1(n340), .IN2(\ram[143][2] ), .IN3(n337), .IN4(
        \ram[144][2] ), .Q(n1163) );
  AOI221X1 U2953 ( .IN1(n373), .IN2(\ram[132][2] ), .IN3(n376), .IN4(
        \ram[131][2] ), .IN5(n1164), .QN(n1161) );
  AO22X1 U2954 ( .IN1(n364), .IN2(\ram[135][2] ), .IN3(n361), .IN4(
        \ram[136][2] ), .Q(n1164) );
  AOI221X1 U2955 ( .IN1(n301), .IN2(\ram[156][2] ), .IN3(n304), .IN4(
        \ram[155][2] ), .IN5(n1165), .QN(n1160) );
  AO22X1 U2956 ( .IN1(n292), .IN2(\ram[159][2] ), .IN3(n289), .IN4(
        \ram[160][2] ), .Q(n1165) );
  AOI221X1 U2957 ( .IN1(n325), .IN2(\ram[148][2] ), .IN3(n328), .IN4(
        \ram[147][2] ), .IN5(n1166), .QN(n1159) );
  AO22X1 U2958 ( .IN1(n316), .IN2(\ram[151][2] ), .IN3(n313), .IN4(
        \ram[152][2] ), .Q(n1166) );
  NAND4X0 U2959 ( .IN1(n1167), .IN2(n1168), .IN3(n1169), .IN4(n1170), .QN(
        n1148) );
  AOI221X1 U2960 ( .IN1(n61), .IN2(\ram[236][2] ), .IN3(n64), .IN4(
        \ram[235][2] ), .IN5(n1171), .QN(n1170) );
  AO22X1 U2961 ( .IN1(n58), .IN2(\ram[237][2] ), .IN3(n55), .IN4(\ram[238][2] ), .Q(n1171) );
  AOI221X1 U2962 ( .IN1(n85), .IN2(\ram[228][2] ), .IN3(n88), .IN4(
        \ram[227][2] ), .IN5(n1172), .QN(n1169) );
  AO22X1 U2963 ( .IN1(n76), .IN2(\ram[231][2] ), .IN3(n73), .IN4(\ram[232][2] ), .Q(n1172) );
  AOI221X1 U2964 ( .IN1(n19), .IN2(\ram[250][2] ), .IN3(n22), .IN4(
        \ram[249][2] ), .IN5(n1173), .QN(n1168) );
  AO22X1 U2965 ( .IN1(n10), .IN2(\ram[253][2] ), .IN3(n7), .IN4(\ram[254][2] ), 
        .Q(n1173) );
  AOI221X1 U2966 ( .IN1(n37), .IN2(\ram[244][2] ), .IN3(n40), .IN4(
        \ram[243][2] ), .IN5(n1174), .QN(n1167) );
  AO22X1 U2967 ( .IN1(n28), .IN2(\ram[247][2] ), .IN3(n25), .IN4(\ram[248][2] ), .Q(n1174) );
  NAND4X0 U2968 ( .IN1(n1175), .IN2(n1176), .IN3(n1177), .IN4(n1178), .QN(
        n1147) );
  AOI221X1 U2969 ( .IN1(n157), .IN2(\ram[204][2] ), .IN3(n160), .IN4(
        \ram[203][2] ), .IN5(n1179), .QN(n1178) );
  AO22X1 U2970 ( .IN1(n148), .IN2(\ram[207][2] ), .IN3(n145), .IN4(
        \ram[208][2] ), .Q(n1179) );
  AOI221X1 U2971 ( .IN1(n181), .IN2(\ram[196][2] ), .IN3(n184), .IN4(
        \ram[195][2] ), .IN5(n1180), .QN(n1177) );
  AO22X1 U2972 ( .IN1(n172), .IN2(\ram[199][2] ), .IN3(n169), .IN4(
        \ram[200][2] ), .Q(n1180) );
  AOI221X1 U2973 ( .IN1(n109), .IN2(\ram[220][2] ), .IN3(n112), .IN4(
        \ram[219][2] ), .IN5(n1181), .QN(n1176) );
  AO22X1 U2974 ( .IN1(n100), .IN2(\ram[223][2] ), .IN3(n97), .IN4(
        \ram[224][2] ), .Q(n1181) );
  AOI221X1 U2975 ( .IN1(n133), .IN2(\ram[212][2] ), .IN3(n136), .IN4(
        \ram[211][2] ), .IN5(n1182), .QN(n1175) );
  AO22X1 U2976 ( .IN1(n124), .IN2(\ram[215][2] ), .IN3(n121), .IN4(
        \ram[216][2] ), .Q(n1182) );
  NAND4X0 U2978 ( .IN1(n1187), .IN2(n1188), .IN3(n1189), .IN4(n1190), .QN(
        n1186) );
  AOI221X1 U2979 ( .IN1(n637), .IN2(\ram[44][2] ), .IN3(n640), .IN4(
        \ram[43][2] ), .IN5(n1191), .QN(n1190) );
  AO22X1 U2980 ( .IN1(n628), .IN2(\ram[47][2] ), .IN3(n625), .IN4(\ram[48][2] ), .Q(n1191) );
  AOI221X1 U2981 ( .IN1(n661), .IN2(\ram[36][2] ), .IN3(n664), .IN4(
        \ram[35][2] ), .IN5(n1192), .QN(n1189) );
  AO22X1 U2982 ( .IN1(n652), .IN2(\ram[39][2] ), .IN3(n649), .IN4(\ram[40][2] ), .Q(n1192) );
  AOI221X1 U2983 ( .IN1(n589), .IN2(\ram[60][2] ), .IN3(n592), .IN4(
        \ram[59][2] ), .IN5(n1193), .QN(n1188) );
  AO22X1 U2984 ( .IN1(n580), .IN2(\ram[63][2] ), .IN3(n577), .IN4(\ram[64][2] ), .Q(n1193) );
  AOI221X1 U2985 ( .IN1(n613), .IN2(\ram[52][2] ), .IN3(n616), .IN4(
        \ram[51][2] ), .IN5(n1194), .QN(n1187) );
  AO22X1 U2986 ( .IN1(n604), .IN2(\ram[55][2] ), .IN3(n601), .IN4(\ram[56][2] ), .Q(n1194) );
  NAND4X0 U2987 ( .IN1(n1195), .IN2(n1196), .IN3(n1197), .IN4(n1198), .QN(
        n1185) );
  AOI221X1 U2988 ( .IN1(n733), .IN2(\ram[12][2] ), .IN3(n736), .IN4(
        \ram[11][2] ), .IN5(n1199), .QN(n1198) );
  AO22X1 U2989 ( .IN1(n724), .IN2(\ram[15][2] ), .IN3(n721), .IN4(\ram[16][2] ), .Q(n1199) );
  AOI221X1 U2990 ( .IN1(n757), .IN2(\ram[4][2] ), .IN3(n760), .IN4(\ram[3][2] ), .IN5(n1200), .QN(n1197) );
  AO22X1 U2991 ( .IN1(n748), .IN2(\ram[7][2] ), .IN3(n745), .IN4(\ram[8][2] ), 
        .Q(n1200) );
  AOI221X1 U2992 ( .IN1(n685), .IN2(\ram[28][2] ), .IN3(n688), .IN4(
        \ram[27][2] ), .IN5(n1201), .QN(n1196) );
  AO22X1 U2993 ( .IN1(n676), .IN2(\ram[31][2] ), .IN3(n673), .IN4(\ram[32][2] ), .Q(n1201) );
  AOI221X1 U2994 ( .IN1(n709), .IN2(\ram[20][2] ), .IN3(n712), .IN4(
        \ram[19][2] ), .IN5(n1202), .QN(n1195) );
  AO22X1 U2995 ( .IN1(n700), .IN2(\ram[23][2] ), .IN3(n697), .IN4(\ram[24][2] ), .Q(n1202) );
  NAND4X0 U2996 ( .IN1(n1203), .IN2(n1204), .IN3(n1205), .IN4(n1206), .QN(
        n1184) );
  AOI221X1 U2997 ( .IN1(n445), .IN2(\ram[108][2] ), .IN3(n448), .IN4(
        \ram[107][2] ), .IN5(n1207), .QN(n1206) );
  AO22X1 U2998 ( .IN1(n436), .IN2(\ram[111][2] ), .IN3(n433), .IN4(
        \ram[112][2] ), .Q(n1207) );
  AOI221X1 U2999 ( .IN1(n469), .IN2(\ram[100][2] ), .IN3(n472), .IN4(
        \ram[99][2] ), .IN5(n1208), .QN(n1205) );
  AO22X1 U3000 ( .IN1(n460), .IN2(\ram[103][2] ), .IN3(n457), .IN4(
        \ram[104][2] ), .Q(n1208) );
  AOI221X1 U3001 ( .IN1(n397), .IN2(\ram[124][2] ), .IN3(n400), .IN4(
        \ram[123][2] ), .IN5(n1209), .QN(n1204) );
  AO22X1 U3002 ( .IN1(n388), .IN2(\ram[127][2] ), .IN3(n385), .IN4(
        \ram[128][2] ), .Q(n1209) );
  AOI221X1 U3003 ( .IN1(n421), .IN2(\ram[116][2] ), .IN3(n424), .IN4(
        \ram[115][2] ), .IN5(n1210), .QN(n1203) );
  AO22X1 U3004 ( .IN1(n412), .IN2(\ram[119][2] ), .IN3(n409), .IN4(
        \ram[120][2] ), .Q(n1210) );
  NAND4X0 U3005 ( .IN1(n1211), .IN2(n1212), .IN3(n1213), .IN4(n1214), .QN(
        n1183) );
  AOI221X1 U3006 ( .IN1(n541), .IN2(\ram[76][2] ), .IN3(n544), .IN4(
        \ram[75][2] ), .IN5(n1215), .QN(n1214) );
  AO22X1 U3007 ( .IN1(n532), .IN2(\ram[79][2] ), .IN3(n529), .IN4(\ram[80][2] ), .Q(n1215) );
  AOI221X1 U3008 ( .IN1(n565), .IN2(\ram[68][2] ), .IN3(n568), .IN4(
        \ram[67][2] ), .IN5(n1216), .QN(n1213) );
  AO22X1 U3009 ( .IN1(n556), .IN2(\ram[71][2] ), .IN3(n553), .IN4(\ram[72][2] ), .Q(n1216) );
  AOI221X1 U3010 ( .IN1(n493), .IN2(\ram[92][2] ), .IN3(n496), .IN4(
        \ram[91][2] ), .IN5(n1217), .QN(n1212) );
  AO22X1 U3011 ( .IN1(n484), .IN2(\ram[95][2] ), .IN3(n481), .IN4(\ram[96][2] ), .Q(n1217) );
  AOI221X1 U3012 ( .IN1(n517), .IN2(\ram[84][2] ), .IN3(n520), .IN4(
        \ram[83][2] ), .IN5(n1218), .QN(n1211) );
  AO22X1 U3013 ( .IN1(n508), .IN2(\ram[87][2] ), .IN3(n505), .IN4(\ram[88][2] ), .Q(n1218) );
  AO22X1 U3014 ( .IN1(n771), .IN2(dataout[3]), .IN3(n4174), .IN4(n1219), .Q(
        n2023) );
  NAND4X0 U3015 ( .IN1(n1220), .IN2(n1221), .IN3(n1222), .IN4(n1223), .QN(
        n1219) );
  NAND4X0 U3017 ( .IN1(n1228), .IN2(n1229), .IN3(n1230), .IN4(n1231), .QN(
        n1227) );
  AOI221X1 U3018 ( .IN1(n259), .IN2(\ram[170][3] ), .IN3(n262), .IN4(
        \ram[169][3] ), .IN5(n1232), .QN(n1231) );
  AO22X1 U3019 ( .IN1(n250), .IN2(\ram[173][3] ), .IN3(n247), .IN4(
        \ram[174][3] ), .Q(n1232) );
  AOI221X1 U3020 ( .IN1(n283), .IN2(\ram[162][3] ), .IN3(n286), .IN4(
        \ram[161][3] ), .IN5(n1233), .QN(n1230) );
  AO22X1 U3021 ( .IN1(n274), .IN2(\ram[165][3] ), .IN3(n271), .IN4(
        \ram[166][3] ), .Q(n1233) );
  AOI221X1 U3022 ( .IN1(n211), .IN2(\ram[186][3] ), .IN3(n214), .IN4(
        \ram[185][3] ), .IN5(n1234), .QN(n1229) );
  AO22X1 U3023 ( .IN1(n196), .IN2(\ram[191][3] ), .IN3(n193), .IN4(
        \ram[192][3] ), .Q(n1234) );
  AOI221X1 U3024 ( .IN1(n235), .IN2(\ram[178][3] ), .IN3(n238), .IN4(
        \ram[177][3] ), .IN5(n1235), .QN(n1228) );
  AO22X1 U3025 ( .IN1(n226), .IN2(\ram[181][3] ), .IN3(n223), .IN4(
        \ram[182][3] ), .Q(n1235) );
  NAND4X0 U3026 ( .IN1(n1236), .IN2(n1237), .IN3(n1238), .IN4(n1239), .QN(
        n1226) );
  AOI221X1 U3027 ( .IN1(n355), .IN2(\ram[138][3] ), .IN3(n358), .IN4(
        \ram[137][3] ), .IN5(n1240), .QN(n1239) );
  AO22X1 U3028 ( .IN1(n346), .IN2(\ram[141][3] ), .IN3(n343), .IN4(
        \ram[142][3] ), .Q(n1240) );
  AOI221X1 U3029 ( .IN1(n379), .IN2(\ram[130][3] ), .IN3(n382), .IN4(
        \ram[129][3] ), .IN5(n1241), .QN(n1238) );
  AO22X1 U3030 ( .IN1(n370), .IN2(\ram[133][3] ), .IN3(n367), .IN4(
        \ram[134][3] ), .Q(n1241) );
  AOI221X1 U3031 ( .IN1(n307), .IN2(\ram[154][3] ), .IN3(n310), .IN4(
        \ram[153][3] ), .IN5(n1242), .QN(n1237) );
  AO22X1 U3032 ( .IN1(n298), .IN2(\ram[157][3] ), .IN3(n295), .IN4(
        \ram[158][3] ), .Q(n1242) );
  AOI221X1 U3033 ( .IN1(n331), .IN2(\ram[146][3] ), .IN3(n334), .IN4(
        \ram[145][3] ), .IN5(n1243), .QN(n1236) );
  AO22X1 U3034 ( .IN1(n322), .IN2(\ram[149][3] ), .IN3(n319), .IN4(
        \ram[150][3] ), .Q(n1243) );
  NAND4X0 U3035 ( .IN1(n1244), .IN2(n1245), .IN3(n1246), .IN4(n1247), .QN(
        n1225) );
  AOI221X1 U3036 ( .IN1(n70), .IN2(\ram[233][3] ), .IN3(n49), .IN4(
        \ram[240][3] ), .IN5(n1248), .QN(n1247) );
  AO22X1 U3037 ( .IN1(n139), .IN2(\ram[210][3] ), .IN3(n52), .IN4(
        \ram[239][3] ), .Q(n1248) );
  AOI221X1 U3038 ( .IN1(n94), .IN2(\ram[225][3] ), .IN3(n79), .IN4(
        \ram[230][3] ), .IN5(n1249), .QN(n1246) );
  AO22X1 U3039 ( .IN1(n67), .IN2(\ram[234][3] ), .IN3(n82), .IN4(\ram[229][3] ), .Q(n1249) );
  AOI221X1 U3040 ( .IN1(n13), .IN2(\ram[252][3] ), .IN3(n16), .IN4(
        \ram[251][3] ), .IN5(n1250), .QN(n1245) );
  AO22X1 U3041 ( .IN1(n91), .IN2(\ram[226][3] ), .IN3(n3), .IN4(\ram[255][3] ), 
        .Q(n1250) );
  AOI221X1 U3042 ( .IN1(n43), .IN2(\ram[242][3] ), .IN3(n46), .IN4(
        \ram[241][3] ), .IN5(n1251), .QN(n1244) );
  AO22X1 U3043 ( .IN1(n34), .IN2(\ram[245][3] ), .IN3(n31), .IN4(\ram[246][3] ), .Q(n1251) );
  NAND4X0 U3044 ( .IN1(n1252), .IN2(n1253), .IN3(n1254), .IN4(n1255), .QN(
        n1224) );
  AOI221X1 U3045 ( .IN1(n166), .IN2(\ram[201][3] ), .IN3(n151), .IN4(
        \ram[206][3] ), .IN5(n1256), .QN(n1255) );
  AO22X1 U3046 ( .IN1(n769), .IN2(\ram[0][3] ), .IN3(n154), .IN4(\ram[205][3] ), .Q(n1256) );
  AOI221X1 U3047 ( .IN1(n190), .IN2(\ram[193][3] ), .IN3(n175), .IN4(
        \ram[198][3] ), .IN5(n1257), .QN(n1254) );
  AO22X1 U3048 ( .IN1(n163), .IN2(\ram[202][3] ), .IN3(n178), .IN4(
        \ram[197][3] ), .Q(n1257) );
  AOI221X1 U3049 ( .IN1(n106), .IN2(\ram[221][3] ), .IN3(n187), .IN4(
        \ram[194][3] ), .IN5(n1258), .QN(n1253) );
  AO22X1 U3050 ( .IN1(n103), .IN2(\ram[222][3] ), .IN3(n118), .IN4(
        \ram[217][3] ), .Q(n1258) );
  AOI221X1 U3051 ( .IN1(n142), .IN2(\ram[209][3] ), .IN3(n127), .IN4(
        \ram[214][3] ), .IN5(n1259), .QN(n1252) );
  AO22X1 U3052 ( .IN1(n115), .IN2(\ram[218][3] ), .IN3(n130), .IN4(
        \ram[213][3] ), .Q(n1259) );
  NAND4X0 U3054 ( .IN1(n1264), .IN2(n1265), .IN3(n1266), .IN4(n1267), .QN(
        n1263) );
  AOI221X1 U3055 ( .IN1(n643), .IN2(\ram[42][3] ), .IN3(n646), .IN4(
        \ram[41][3] ), .IN5(n1268), .QN(n1267) );
  AO22X1 U3056 ( .IN1(n634), .IN2(\ram[45][3] ), .IN3(n631), .IN4(\ram[46][3] ), .Q(n1268) );
  AOI221X1 U3057 ( .IN1(n667), .IN2(\ram[34][3] ), .IN3(n670), .IN4(
        \ram[33][3] ), .IN5(n1269), .QN(n1266) );
  AO22X1 U3058 ( .IN1(n658), .IN2(\ram[37][3] ), .IN3(n655), .IN4(\ram[38][3] ), .Q(n1269) );
  AOI221X1 U3059 ( .IN1(n595), .IN2(\ram[58][3] ), .IN3(n598), .IN4(
        \ram[57][3] ), .IN5(n1270), .QN(n1265) );
  AO22X1 U3060 ( .IN1(n586), .IN2(\ram[61][3] ), .IN3(n583), .IN4(\ram[62][3] ), .Q(n1270) );
  AOI221X1 U3061 ( .IN1(n619), .IN2(\ram[50][3] ), .IN3(n622), .IN4(
        \ram[49][3] ), .IN5(n1271), .QN(n1264) );
  AO22X1 U3062 ( .IN1(n610), .IN2(\ram[53][3] ), .IN3(n607), .IN4(\ram[54][3] ), .Q(n1271) );
  NAND4X0 U3063 ( .IN1(n1272), .IN2(n1273), .IN3(n1274), .IN4(n1275), .QN(
        n1262) );
  AOI221X1 U3064 ( .IN1(n739), .IN2(\ram[10][3] ), .IN3(n742), .IN4(
        \ram[9][3] ), .IN5(n1276), .QN(n1275) );
  AO22X1 U3065 ( .IN1(n730), .IN2(\ram[13][3] ), .IN3(n727), .IN4(\ram[14][3] ), .Q(n1276) );
  AOI221X1 U3066 ( .IN1(n763), .IN2(\ram[2][3] ), .IN3(n766), .IN4(\ram[1][3] ), .IN5(n1277), .QN(n1274) );
  AO22X1 U3067 ( .IN1(n754), .IN2(\ram[5][3] ), .IN3(n751), .IN4(\ram[6][3] ), 
        .Q(n1277) );
  AOI221X1 U3068 ( .IN1(n691), .IN2(\ram[26][3] ), .IN3(n694), .IN4(
        \ram[25][3] ), .IN5(n1278), .QN(n1273) );
  AO22X1 U3069 ( .IN1(n682), .IN2(\ram[29][3] ), .IN3(n679), .IN4(\ram[30][3] ), .Q(n1278) );
  AOI221X1 U3070 ( .IN1(n715), .IN2(\ram[18][3] ), .IN3(n718), .IN4(
        \ram[17][3] ), .IN5(n1279), .QN(n1272) );
  AO22X1 U3071 ( .IN1(n706), .IN2(\ram[21][3] ), .IN3(n703), .IN4(\ram[22][3] ), .Q(n1279) );
  NAND4X0 U3072 ( .IN1(n1280), .IN2(n1281), .IN3(n1282), .IN4(n1283), .QN(
        n1261) );
  AOI221X1 U3073 ( .IN1(n451), .IN2(\ram[106][3] ), .IN3(n454), .IN4(
        \ram[105][3] ), .IN5(n1284), .QN(n1283) );
  AO22X1 U3074 ( .IN1(n442), .IN2(\ram[109][3] ), .IN3(n439), .IN4(
        \ram[110][3] ), .Q(n1284) );
  AOI221X1 U3075 ( .IN1(n475), .IN2(\ram[98][3] ), .IN3(n478), .IN4(
        \ram[97][3] ), .IN5(n1285), .QN(n1282) );
  AO22X1 U3076 ( .IN1(n466), .IN2(\ram[101][3] ), .IN3(n463), .IN4(
        \ram[102][3] ), .Q(n1285) );
  AOI221X1 U3077 ( .IN1(n403), .IN2(\ram[122][3] ), .IN3(n406), .IN4(
        \ram[121][3] ), .IN5(n1286), .QN(n1281) );
  AO22X1 U3078 ( .IN1(n394), .IN2(\ram[125][3] ), .IN3(n391), .IN4(
        \ram[126][3] ), .Q(n1286) );
  AOI221X1 U3079 ( .IN1(n427), .IN2(\ram[114][3] ), .IN3(n430), .IN4(
        \ram[113][3] ), .IN5(n1287), .QN(n1280) );
  AO22X1 U3080 ( .IN1(n418), .IN2(\ram[117][3] ), .IN3(n415), .IN4(
        \ram[118][3] ), .Q(n1287) );
  NAND4X0 U3081 ( .IN1(n1288), .IN2(n1289), .IN3(n1290), .IN4(n1291), .QN(
        n1260) );
  AOI221X1 U3082 ( .IN1(n547), .IN2(\ram[74][3] ), .IN3(n550), .IN4(
        \ram[73][3] ), .IN5(n1292), .QN(n1291) );
  AO22X1 U3083 ( .IN1(n538), .IN2(\ram[77][3] ), .IN3(n535), .IN4(\ram[78][3] ), .Q(n1292) );
  AOI221X1 U3084 ( .IN1(n571), .IN2(\ram[66][3] ), .IN3(n574), .IN4(
        \ram[65][3] ), .IN5(n1293), .QN(n1290) );
  AO22X1 U3085 ( .IN1(n562), .IN2(\ram[69][3] ), .IN3(n559), .IN4(\ram[70][3] ), .Q(n1293) );
  AOI221X1 U3086 ( .IN1(n499), .IN2(\ram[90][3] ), .IN3(n502), .IN4(
        \ram[89][3] ), .IN5(n1294), .QN(n1289) );
  AO22X1 U3087 ( .IN1(n490), .IN2(\ram[93][3] ), .IN3(n487), .IN4(\ram[94][3] ), .Q(n1294) );
  AOI221X1 U3088 ( .IN1(n523), .IN2(\ram[82][3] ), .IN3(n526), .IN4(
        \ram[81][3] ), .IN5(n1295), .QN(n1288) );
  AO22X1 U3089 ( .IN1(n514), .IN2(\ram[85][3] ), .IN3(n511), .IN4(\ram[86][3] ), .Q(n1295) );
  NAND4X0 U3091 ( .IN1(n1300), .IN2(n1301), .IN3(n1302), .IN4(n1303), .QN(
        n1299) );
  AOI221X1 U3092 ( .IN1(n253), .IN2(\ram[172][3] ), .IN3(n256), .IN4(
        \ram[171][3] ), .IN5(n1304), .QN(n1303) );
  AO22X1 U3093 ( .IN1(n244), .IN2(\ram[175][3] ), .IN3(n241), .IN4(
        \ram[176][3] ), .Q(n1304) );
  AOI221X1 U3094 ( .IN1(n277), .IN2(\ram[164][3] ), .IN3(n280), .IN4(
        \ram[163][3] ), .IN5(n1305), .QN(n1302) );
  AO22X1 U3095 ( .IN1(n268), .IN2(\ram[167][3] ), .IN3(n265), .IN4(
        \ram[168][3] ), .Q(n1305) );
  AOI221X1 U3096 ( .IN1(n205), .IN2(\ram[188][3] ), .IN3(n208), .IN4(
        \ram[187][3] ), .IN5(n1306), .QN(n1301) );
  AO22X1 U3097 ( .IN1(n202), .IN2(\ram[189][3] ), .IN3(n199), .IN4(
        \ram[190][3] ), .Q(n1306) );
  AOI221X1 U3098 ( .IN1(n229), .IN2(\ram[180][3] ), .IN3(n232), .IN4(
        \ram[179][3] ), .IN5(n1307), .QN(n1300) );
  AO22X1 U3099 ( .IN1(n220), .IN2(\ram[183][3] ), .IN3(n217), .IN4(
        \ram[184][3] ), .Q(n1307) );
  NAND4X0 U3100 ( .IN1(n1308), .IN2(n1309), .IN3(n1310), .IN4(n1311), .QN(
        n1298) );
  AOI221X1 U3101 ( .IN1(n349), .IN2(\ram[140][3] ), .IN3(n352), .IN4(
        \ram[139][3] ), .IN5(n1312), .QN(n1311) );
  AO22X1 U3102 ( .IN1(n340), .IN2(\ram[143][3] ), .IN3(n337), .IN4(
        \ram[144][3] ), .Q(n1312) );
  AOI221X1 U3103 ( .IN1(n373), .IN2(\ram[132][3] ), .IN3(n376), .IN4(
        \ram[131][3] ), .IN5(n1313), .QN(n1310) );
  AO22X1 U3104 ( .IN1(n364), .IN2(\ram[135][3] ), .IN3(n361), .IN4(
        \ram[136][3] ), .Q(n1313) );
  AOI221X1 U3105 ( .IN1(n301), .IN2(\ram[156][3] ), .IN3(n304), .IN4(
        \ram[155][3] ), .IN5(n1314), .QN(n1309) );
  AO22X1 U3106 ( .IN1(n292), .IN2(\ram[159][3] ), .IN3(n289), .IN4(
        \ram[160][3] ), .Q(n1314) );
  AOI221X1 U3107 ( .IN1(n325), .IN2(\ram[148][3] ), .IN3(n328), .IN4(
        \ram[147][3] ), .IN5(n1315), .QN(n1308) );
  AO22X1 U3108 ( .IN1(n316), .IN2(\ram[151][3] ), .IN3(n313), .IN4(
        \ram[152][3] ), .Q(n1315) );
  NAND4X0 U3109 ( .IN1(n1316), .IN2(n1317), .IN3(n1318), .IN4(n1319), .QN(
        n1297) );
  AOI221X1 U3110 ( .IN1(n61), .IN2(\ram[236][3] ), .IN3(n64), .IN4(
        \ram[235][3] ), .IN5(n1320), .QN(n1319) );
  AO22X1 U3111 ( .IN1(n58), .IN2(\ram[237][3] ), .IN3(n55), .IN4(\ram[238][3] ), .Q(n1320) );
  AOI221X1 U3112 ( .IN1(n85), .IN2(\ram[228][3] ), .IN3(n88), .IN4(
        \ram[227][3] ), .IN5(n1321), .QN(n1318) );
  AO22X1 U3113 ( .IN1(n76), .IN2(\ram[231][3] ), .IN3(n73), .IN4(\ram[232][3] ), .Q(n1321) );
  AOI221X1 U3114 ( .IN1(n19), .IN2(\ram[250][3] ), .IN3(n22), .IN4(
        \ram[249][3] ), .IN5(n1322), .QN(n1317) );
  AO22X1 U3115 ( .IN1(n10), .IN2(\ram[253][3] ), .IN3(n7), .IN4(\ram[254][3] ), 
        .Q(n1322) );
  AOI221X1 U3116 ( .IN1(n37), .IN2(\ram[244][3] ), .IN3(n40), .IN4(
        \ram[243][3] ), .IN5(n1323), .QN(n1316) );
  AO22X1 U3117 ( .IN1(n28), .IN2(\ram[247][3] ), .IN3(n25), .IN4(\ram[248][3] ), .Q(n1323) );
  NAND4X0 U3118 ( .IN1(n1324), .IN2(n1325), .IN3(n1326), .IN4(n1327), .QN(
        n1296) );
  AOI221X1 U3119 ( .IN1(n157), .IN2(\ram[204][3] ), .IN3(n160), .IN4(
        \ram[203][3] ), .IN5(n1328), .QN(n1327) );
  AO22X1 U3120 ( .IN1(n148), .IN2(\ram[207][3] ), .IN3(n145), .IN4(
        \ram[208][3] ), .Q(n1328) );
  AOI221X1 U3121 ( .IN1(n181), .IN2(\ram[196][3] ), .IN3(n184), .IN4(
        \ram[195][3] ), .IN5(n1329), .QN(n1326) );
  AO22X1 U3122 ( .IN1(n172), .IN2(\ram[199][3] ), .IN3(n169), .IN4(
        \ram[200][3] ), .Q(n1329) );
  AOI221X1 U3123 ( .IN1(n109), .IN2(\ram[220][3] ), .IN3(n112), .IN4(
        \ram[219][3] ), .IN5(n1330), .QN(n1325) );
  AO22X1 U3124 ( .IN1(n100), .IN2(\ram[223][3] ), .IN3(n97), .IN4(
        \ram[224][3] ), .Q(n1330) );
  AOI221X1 U3125 ( .IN1(n133), .IN2(\ram[212][3] ), .IN3(n136), .IN4(
        \ram[211][3] ), .IN5(n1331), .QN(n1324) );
  AO22X1 U3126 ( .IN1(n124), .IN2(\ram[215][3] ), .IN3(n121), .IN4(
        \ram[216][3] ), .Q(n1331) );
  NAND4X0 U3128 ( .IN1(n1336), .IN2(n1337), .IN3(n1338), .IN4(n1339), .QN(
        n1335) );
  AOI221X1 U3129 ( .IN1(n637), .IN2(\ram[44][3] ), .IN3(n640), .IN4(
        \ram[43][3] ), .IN5(n1340), .QN(n1339) );
  AO22X1 U3130 ( .IN1(n628), .IN2(\ram[47][3] ), .IN3(n625), .IN4(\ram[48][3] ), .Q(n1340) );
  AOI221X1 U3131 ( .IN1(n661), .IN2(\ram[36][3] ), .IN3(n664), .IN4(
        \ram[35][3] ), .IN5(n1341), .QN(n1338) );
  AO22X1 U3132 ( .IN1(n652), .IN2(\ram[39][3] ), .IN3(n649), .IN4(\ram[40][3] ), .Q(n1341) );
  AOI221X1 U3133 ( .IN1(n589), .IN2(\ram[60][3] ), .IN3(n592), .IN4(
        \ram[59][3] ), .IN5(n1342), .QN(n1337) );
  AO22X1 U3134 ( .IN1(n580), .IN2(\ram[63][3] ), .IN3(n577), .IN4(\ram[64][3] ), .Q(n1342) );
  AOI221X1 U3135 ( .IN1(n613), .IN2(\ram[52][3] ), .IN3(n616), .IN4(
        \ram[51][3] ), .IN5(n1343), .QN(n1336) );
  AO22X1 U3136 ( .IN1(n604), .IN2(\ram[55][3] ), .IN3(n601), .IN4(\ram[56][3] ), .Q(n1343) );
  NAND4X0 U3137 ( .IN1(n1344), .IN2(n1345), .IN3(n1346), .IN4(n1347), .QN(
        n1334) );
  AOI221X1 U3138 ( .IN1(n733), .IN2(\ram[12][3] ), .IN3(n736), .IN4(
        \ram[11][3] ), .IN5(n1348), .QN(n1347) );
  AO22X1 U3139 ( .IN1(n724), .IN2(\ram[15][3] ), .IN3(n721), .IN4(\ram[16][3] ), .Q(n1348) );
  AOI221X1 U3140 ( .IN1(n757), .IN2(\ram[4][3] ), .IN3(n760), .IN4(\ram[3][3] ), .IN5(n1349), .QN(n1346) );
  AO22X1 U3141 ( .IN1(n748), .IN2(\ram[7][3] ), .IN3(n745), .IN4(\ram[8][3] ), 
        .Q(n1349) );
  AOI221X1 U3142 ( .IN1(n685), .IN2(\ram[28][3] ), .IN3(n688), .IN4(
        \ram[27][3] ), .IN5(n1350), .QN(n1345) );
  AO22X1 U3143 ( .IN1(n676), .IN2(\ram[31][3] ), .IN3(n673), .IN4(\ram[32][3] ), .Q(n1350) );
  AOI221X1 U3144 ( .IN1(n709), .IN2(\ram[20][3] ), .IN3(n712), .IN4(
        \ram[19][3] ), .IN5(n1351), .QN(n1344) );
  AO22X1 U3145 ( .IN1(n700), .IN2(\ram[23][3] ), .IN3(n697), .IN4(\ram[24][3] ), .Q(n1351) );
  NAND4X0 U3146 ( .IN1(n1352), .IN2(n1353), .IN3(n1354), .IN4(n1355), .QN(
        n1333) );
  AOI221X1 U3147 ( .IN1(n445), .IN2(\ram[108][3] ), .IN3(n448), .IN4(
        \ram[107][3] ), .IN5(n1356), .QN(n1355) );
  AO22X1 U3148 ( .IN1(n436), .IN2(\ram[111][3] ), .IN3(n433), .IN4(
        \ram[112][3] ), .Q(n1356) );
  AOI221X1 U3149 ( .IN1(n469), .IN2(\ram[100][3] ), .IN3(n472), .IN4(
        \ram[99][3] ), .IN5(n1357), .QN(n1354) );
  AO22X1 U3150 ( .IN1(n460), .IN2(\ram[103][3] ), .IN3(n457), .IN4(
        \ram[104][3] ), .Q(n1357) );
  AOI221X1 U3151 ( .IN1(n397), .IN2(\ram[124][3] ), .IN3(n400), .IN4(
        \ram[123][3] ), .IN5(n1358), .QN(n1353) );
  AO22X1 U3152 ( .IN1(n388), .IN2(\ram[127][3] ), .IN3(n385), .IN4(
        \ram[128][3] ), .Q(n1358) );
  AOI221X1 U3153 ( .IN1(n421), .IN2(\ram[116][3] ), .IN3(n424), .IN4(
        \ram[115][3] ), .IN5(n1359), .QN(n1352) );
  AO22X1 U3154 ( .IN1(n412), .IN2(\ram[119][3] ), .IN3(n409), .IN4(
        \ram[120][3] ), .Q(n1359) );
  NAND4X0 U3155 ( .IN1(n1360), .IN2(n1361), .IN3(n1362), .IN4(n1363), .QN(
        n1332) );
  AOI221X1 U3156 ( .IN1(n541), .IN2(\ram[76][3] ), .IN3(n544), .IN4(
        \ram[75][3] ), .IN5(n1364), .QN(n1363) );
  AO22X1 U3157 ( .IN1(n532), .IN2(\ram[79][3] ), .IN3(n529), .IN4(\ram[80][3] ), .Q(n1364) );
  AOI221X1 U3158 ( .IN1(n565), .IN2(\ram[68][3] ), .IN3(n568), .IN4(
        \ram[67][3] ), .IN5(n1365), .QN(n1362) );
  AO22X1 U3159 ( .IN1(n556), .IN2(\ram[71][3] ), .IN3(n553), .IN4(\ram[72][3] ), .Q(n1365) );
  AOI221X1 U3160 ( .IN1(n493), .IN2(\ram[92][3] ), .IN3(n496), .IN4(
        \ram[91][3] ), .IN5(n1366), .QN(n1361) );
  AO22X1 U3161 ( .IN1(n484), .IN2(\ram[95][3] ), .IN3(n481), .IN4(\ram[96][3] ), .Q(n1366) );
  AOI221X1 U3162 ( .IN1(n517), .IN2(\ram[84][3] ), .IN3(n520), .IN4(
        \ram[83][3] ), .IN5(n1367), .QN(n1360) );
  AO22X1 U3163 ( .IN1(n508), .IN2(\ram[87][3] ), .IN3(n505), .IN4(\ram[88][3] ), .Q(n1367) );
  AO22X1 U3164 ( .IN1(n771), .IN2(dataout[4]), .IN3(n4174), .IN4(n1368), .Q(
        n2024) );
  NAND4X0 U3165 ( .IN1(n1369), .IN2(n1370), .IN3(n1371), .IN4(n1372), .QN(
        n1368) );
  NAND4X0 U3167 ( .IN1(n1377), .IN2(n1378), .IN3(n1379), .IN4(n1380), .QN(
        n1376) );
  AOI221X1 U3168 ( .IN1(n259), .IN2(\ram[170][4] ), .IN3(n262), .IN4(
        \ram[169][4] ), .IN5(n1381), .QN(n1380) );
  AO22X1 U3169 ( .IN1(n250), .IN2(\ram[173][4] ), .IN3(n247), .IN4(
        \ram[174][4] ), .Q(n1381) );
  AOI221X1 U3170 ( .IN1(n283), .IN2(\ram[162][4] ), .IN3(n286), .IN4(
        \ram[161][4] ), .IN5(n1382), .QN(n1379) );
  AO22X1 U3171 ( .IN1(n274), .IN2(\ram[165][4] ), .IN3(n271), .IN4(
        \ram[166][4] ), .Q(n1382) );
  AOI221X1 U3172 ( .IN1(n211), .IN2(\ram[186][4] ), .IN3(n214), .IN4(
        \ram[185][4] ), .IN5(n1383), .QN(n1378) );
  AO22X1 U3173 ( .IN1(n196), .IN2(\ram[191][4] ), .IN3(n193), .IN4(
        \ram[192][4] ), .Q(n1383) );
  AOI221X1 U3174 ( .IN1(n235), .IN2(\ram[178][4] ), .IN3(n238), .IN4(
        \ram[177][4] ), .IN5(n1384), .QN(n1377) );
  AO22X1 U3175 ( .IN1(n226), .IN2(\ram[181][4] ), .IN3(n223), .IN4(
        \ram[182][4] ), .Q(n1384) );
  NAND4X0 U3176 ( .IN1(n1385), .IN2(n1386), .IN3(n1387), .IN4(n1388), .QN(
        n1375) );
  AOI221X1 U3177 ( .IN1(n355), .IN2(\ram[138][4] ), .IN3(n358), .IN4(
        \ram[137][4] ), .IN5(n1389), .QN(n1388) );
  AO22X1 U3178 ( .IN1(n346), .IN2(\ram[141][4] ), .IN3(n343), .IN4(
        \ram[142][4] ), .Q(n1389) );
  AOI221X1 U3179 ( .IN1(n379), .IN2(\ram[130][4] ), .IN3(n382), .IN4(
        \ram[129][4] ), .IN5(n1390), .QN(n1387) );
  AO22X1 U3180 ( .IN1(n370), .IN2(\ram[133][4] ), .IN3(n367), .IN4(
        \ram[134][4] ), .Q(n1390) );
  AOI221X1 U3181 ( .IN1(n307), .IN2(\ram[154][4] ), .IN3(n310), .IN4(
        \ram[153][4] ), .IN5(n1391), .QN(n1386) );
  AO22X1 U3182 ( .IN1(n298), .IN2(\ram[157][4] ), .IN3(n295), .IN4(
        \ram[158][4] ), .Q(n1391) );
  AOI221X1 U3183 ( .IN1(n331), .IN2(\ram[146][4] ), .IN3(n334), .IN4(
        \ram[145][4] ), .IN5(n1392), .QN(n1385) );
  AO22X1 U3184 ( .IN1(n322), .IN2(\ram[149][4] ), .IN3(n319), .IN4(
        \ram[150][4] ), .Q(n1392) );
  NAND4X0 U3185 ( .IN1(n1393), .IN2(n1394), .IN3(n1395), .IN4(n1396), .QN(
        n1374) );
  AOI221X1 U3186 ( .IN1(n70), .IN2(\ram[233][4] ), .IN3(n49), .IN4(
        \ram[240][4] ), .IN5(n1397), .QN(n1396) );
  AO22X1 U3187 ( .IN1(n139), .IN2(\ram[210][4] ), .IN3(n52), .IN4(
        \ram[239][4] ), .Q(n1397) );
  AOI221X1 U3188 ( .IN1(n94), .IN2(\ram[225][4] ), .IN3(n79), .IN4(
        \ram[230][4] ), .IN5(n1398), .QN(n1395) );
  AO22X1 U3189 ( .IN1(n67), .IN2(\ram[234][4] ), .IN3(n82), .IN4(\ram[229][4] ), .Q(n1398) );
  AOI221X1 U3190 ( .IN1(n13), .IN2(\ram[252][4] ), .IN3(n16), .IN4(
        \ram[251][4] ), .IN5(n1399), .QN(n1394) );
  AO22X1 U3191 ( .IN1(n91), .IN2(\ram[226][4] ), .IN3(n3), .IN4(\ram[255][4] ), 
        .Q(n1399) );
  AOI221X1 U3192 ( .IN1(n43), .IN2(\ram[242][4] ), .IN3(n46), .IN4(
        \ram[241][4] ), .IN5(n1400), .QN(n1393) );
  AO22X1 U3193 ( .IN1(n34), .IN2(\ram[245][4] ), .IN3(n31), .IN4(\ram[246][4] ), .Q(n1400) );
  NAND4X0 U3194 ( .IN1(n1401), .IN2(n1402), .IN3(n1403), .IN4(n1404), .QN(
        n1373) );
  AOI221X1 U3195 ( .IN1(n166), .IN2(\ram[201][4] ), .IN3(n151), .IN4(
        \ram[206][4] ), .IN5(n1405), .QN(n1404) );
  AO22X1 U3196 ( .IN1(n769), .IN2(\ram[0][4] ), .IN3(n154), .IN4(\ram[205][4] ), .Q(n1405) );
  AOI221X1 U3197 ( .IN1(n190), .IN2(\ram[193][4] ), .IN3(n175), .IN4(
        \ram[198][4] ), .IN5(n1406), .QN(n1403) );
  AO22X1 U3198 ( .IN1(n163), .IN2(\ram[202][4] ), .IN3(n178), .IN4(
        \ram[197][4] ), .Q(n1406) );
  AOI221X1 U3199 ( .IN1(n106), .IN2(\ram[221][4] ), .IN3(n187), .IN4(
        \ram[194][4] ), .IN5(n1407), .QN(n1402) );
  AO22X1 U3200 ( .IN1(n103), .IN2(\ram[222][4] ), .IN3(n118), .IN4(
        \ram[217][4] ), .Q(n1407) );
  AOI221X1 U3201 ( .IN1(n142), .IN2(\ram[209][4] ), .IN3(n127), .IN4(
        \ram[214][4] ), .IN5(n1408), .QN(n1401) );
  AO22X1 U3202 ( .IN1(n115), .IN2(\ram[218][4] ), .IN3(n130), .IN4(
        \ram[213][4] ), .Q(n1408) );
  NAND4X0 U3204 ( .IN1(n1413), .IN2(n1414), .IN3(n1415), .IN4(n1416), .QN(
        n1412) );
  AOI221X1 U3205 ( .IN1(n643), .IN2(\ram[42][4] ), .IN3(n646), .IN4(
        \ram[41][4] ), .IN5(n1417), .QN(n1416) );
  AO22X1 U3206 ( .IN1(n634), .IN2(\ram[45][4] ), .IN3(n631), .IN4(\ram[46][4] ), .Q(n1417) );
  AOI221X1 U3207 ( .IN1(n667), .IN2(\ram[34][4] ), .IN3(n670), .IN4(
        \ram[33][4] ), .IN5(n1418), .QN(n1415) );
  AO22X1 U3208 ( .IN1(n658), .IN2(\ram[37][4] ), .IN3(n655), .IN4(\ram[38][4] ), .Q(n1418) );
  AOI221X1 U3209 ( .IN1(n595), .IN2(\ram[58][4] ), .IN3(n598), .IN4(
        \ram[57][4] ), .IN5(n1419), .QN(n1414) );
  AO22X1 U3210 ( .IN1(n586), .IN2(\ram[61][4] ), .IN3(n583), .IN4(\ram[62][4] ), .Q(n1419) );
  AOI221X1 U3211 ( .IN1(n619), .IN2(\ram[50][4] ), .IN3(n622), .IN4(
        \ram[49][4] ), .IN5(n1420), .QN(n1413) );
  AO22X1 U3212 ( .IN1(n610), .IN2(\ram[53][4] ), .IN3(n607), .IN4(\ram[54][4] ), .Q(n1420) );
  NAND4X0 U3213 ( .IN1(n1421), .IN2(n1422), .IN3(n1423), .IN4(n1424), .QN(
        n1411) );
  AOI221X1 U3214 ( .IN1(n739), .IN2(\ram[10][4] ), .IN3(n742), .IN4(
        \ram[9][4] ), .IN5(n1425), .QN(n1424) );
  AO22X1 U3215 ( .IN1(n730), .IN2(\ram[13][4] ), .IN3(n727), .IN4(\ram[14][4] ), .Q(n1425) );
  AOI221X1 U3216 ( .IN1(n763), .IN2(\ram[2][4] ), .IN3(n766), .IN4(\ram[1][4] ), .IN5(n1426), .QN(n1423) );
  AO22X1 U3217 ( .IN1(n754), .IN2(\ram[5][4] ), .IN3(n751), .IN4(\ram[6][4] ), 
        .Q(n1426) );
  AOI221X1 U3218 ( .IN1(n691), .IN2(\ram[26][4] ), .IN3(n694), .IN4(
        \ram[25][4] ), .IN5(n1427), .QN(n1422) );
  AO22X1 U3219 ( .IN1(n682), .IN2(\ram[29][4] ), .IN3(n679), .IN4(\ram[30][4] ), .Q(n1427) );
  AOI221X1 U3220 ( .IN1(n715), .IN2(\ram[18][4] ), .IN3(n718), .IN4(
        \ram[17][4] ), .IN5(n1428), .QN(n1421) );
  AO22X1 U3221 ( .IN1(n706), .IN2(\ram[21][4] ), .IN3(n703), .IN4(\ram[22][4] ), .Q(n1428) );
  NAND4X0 U3222 ( .IN1(n1429), .IN2(n1430), .IN3(n1431), .IN4(n1432), .QN(
        n1410) );
  AOI221X1 U3223 ( .IN1(n451), .IN2(\ram[106][4] ), .IN3(n454), .IN4(
        \ram[105][4] ), .IN5(n1433), .QN(n1432) );
  AO22X1 U3224 ( .IN1(n442), .IN2(\ram[109][4] ), .IN3(n439), .IN4(
        \ram[110][4] ), .Q(n1433) );
  AOI221X1 U3225 ( .IN1(n475), .IN2(\ram[98][4] ), .IN3(n478), .IN4(
        \ram[97][4] ), .IN5(n1434), .QN(n1431) );
  AO22X1 U3226 ( .IN1(n466), .IN2(\ram[101][4] ), .IN3(n463), .IN4(
        \ram[102][4] ), .Q(n1434) );
  AOI221X1 U3227 ( .IN1(n403), .IN2(\ram[122][4] ), .IN3(n406), .IN4(
        \ram[121][4] ), .IN5(n1435), .QN(n1430) );
  AO22X1 U3228 ( .IN1(n394), .IN2(\ram[125][4] ), .IN3(n391), .IN4(
        \ram[126][4] ), .Q(n1435) );
  AOI221X1 U3229 ( .IN1(n427), .IN2(\ram[114][4] ), .IN3(n430), .IN4(
        \ram[113][4] ), .IN5(n1436), .QN(n1429) );
  AO22X1 U3230 ( .IN1(n418), .IN2(\ram[117][4] ), .IN3(n415), .IN4(
        \ram[118][4] ), .Q(n1436) );
  NAND4X0 U3231 ( .IN1(n1437), .IN2(n1438), .IN3(n1439), .IN4(n1440), .QN(
        n1409) );
  AOI221X1 U3232 ( .IN1(n547), .IN2(\ram[74][4] ), .IN3(n550), .IN4(
        \ram[73][4] ), .IN5(n1441), .QN(n1440) );
  AO22X1 U3233 ( .IN1(n538), .IN2(\ram[77][4] ), .IN3(n535), .IN4(\ram[78][4] ), .Q(n1441) );
  AOI221X1 U3234 ( .IN1(n571), .IN2(\ram[66][4] ), .IN3(n574), .IN4(
        \ram[65][4] ), .IN5(n1442), .QN(n1439) );
  AO22X1 U3235 ( .IN1(n562), .IN2(\ram[69][4] ), .IN3(n559), .IN4(\ram[70][4] ), .Q(n1442) );
  AOI221X1 U3236 ( .IN1(n499), .IN2(\ram[90][4] ), .IN3(n502), .IN4(
        \ram[89][4] ), .IN5(n1443), .QN(n1438) );
  AO22X1 U3237 ( .IN1(n490), .IN2(\ram[93][4] ), .IN3(n487), .IN4(\ram[94][4] ), .Q(n1443) );
  AOI221X1 U3238 ( .IN1(n523), .IN2(\ram[82][4] ), .IN3(n526), .IN4(
        \ram[81][4] ), .IN5(n1444), .QN(n1437) );
  AO22X1 U3239 ( .IN1(n514), .IN2(\ram[85][4] ), .IN3(n511), .IN4(\ram[86][4] ), .Q(n1444) );
  NAND4X0 U3241 ( .IN1(n1449), .IN2(n1450), .IN3(n1451), .IN4(n1452), .QN(
        n1448) );
  AOI221X1 U3242 ( .IN1(n253), .IN2(\ram[172][4] ), .IN3(n256), .IN4(
        \ram[171][4] ), .IN5(n1453), .QN(n1452) );
  AO22X1 U3243 ( .IN1(n244), .IN2(\ram[175][4] ), .IN3(n241), .IN4(
        \ram[176][4] ), .Q(n1453) );
  AOI221X1 U3244 ( .IN1(n277), .IN2(\ram[164][4] ), .IN3(n280), .IN4(
        \ram[163][4] ), .IN5(n1454), .QN(n1451) );
  AO22X1 U3245 ( .IN1(n268), .IN2(\ram[167][4] ), .IN3(n265), .IN4(
        \ram[168][4] ), .Q(n1454) );
  AOI221X1 U3246 ( .IN1(n205), .IN2(\ram[188][4] ), .IN3(n208), .IN4(
        \ram[187][4] ), .IN5(n1455), .QN(n1450) );
  AO22X1 U3247 ( .IN1(n202), .IN2(\ram[189][4] ), .IN3(n199), .IN4(
        \ram[190][4] ), .Q(n1455) );
  AOI221X1 U3248 ( .IN1(n229), .IN2(\ram[180][4] ), .IN3(n232), .IN4(
        \ram[179][4] ), .IN5(n1456), .QN(n1449) );
  AO22X1 U3249 ( .IN1(n220), .IN2(\ram[183][4] ), .IN3(n217), .IN4(
        \ram[184][4] ), .Q(n1456) );
  NAND4X0 U3250 ( .IN1(n1457), .IN2(n1458), .IN3(n1459), .IN4(n1460), .QN(
        n1447) );
  AOI221X1 U3251 ( .IN1(n349), .IN2(\ram[140][4] ), .IN3(n352), .IN4(
        \ram[139][4] ), .IN5(n1461), .QN(n1460) );
  AO22X1 U3252 ( .IN1(n340), .IN2(\ram[143][4] ), .IN3(n337), .IN4(
        \ram[144][4] ), .Q(n1461) );
  AOI221X1 U3253 ( .IN1(n373), .IN2(\ram[132][4] ), .IN3(n376), .IN4(
        \ram[131][4] ), .IN5(n1462), .QN(n1459) );
  AO22X1 U3254 ( .IN1(n364), .IN2(\ram[135][4] ), .IN3(n361), .IN4(
        \ram[136][4] ), .Q(n1462) );
  AOI221X1 U3255 ( .IN1(n301), .IN2(\ram[156][4] ), .IN3(n304), .IN4(
        \ram[155][4] ), .IN5(n1463), .QN(n1458) );
  AO22X1 U3256 ( .IN1(n292), .IN2(\ram[159][4] ), .IN3(n289), .IN4(
        \ram[160][4] ), .Q(n1463) );
  AOI221X1 U3257 ( .IN1(n325), .IN2(\ram[148][4] ), .IN3(n328), .IN4(
        \ram[147][4] ), .IN5(n1464), .QN(n1457) );
  AO22X1 U3258 ( .IN1(n316), .IN2(\ram[151][4] ), .IN3(n313), .IN4(
        \ram[152][4] ), .Q(n1464) );
  NAND4X0 U3259 ( .IN1(n1465), .IN2(n1466), .IN3(n1467), .IN4(n1468), .QN(
        n1446) );
  AOI221X1 U3260 ( .IN1(n61), .IN2(\ram[236][4] ), .IN3(n64), .IN4(
        \ram[235][4] ), .IN5(n1469), .QN(n1468) );
  AO22X1 U3261 ( .IN1(n58), .IN2(\ram[237][4] ), .IN3(n55), .IN4(\ram[238][4] ), .Q(n1469) );
  AOI221X1 U3262 ( .IN1(n85), .IN2(\ram[228][4] ), .IN3(n88), .IN4(
        \ram[227][4] ), .IN5(n1470), .QN(n1467) );
  AO22X1 U3263 ( .IN1(n76), .IN2(\ram[231][4] ), .IN3(n73), .IN4(\ram[232][4] ), .Q(n1470) );
  AOI221X1 U3264 ( .IN1(n19), .IN2(\ram[250][4] ), .IN3(n22), .IN4(
        \ram[249][4] ), .IN5(n1471), .QN(n1466) );
  AO22X1 U3265 ( .IN1(n10), .IN2(\ram[253][4] ), .IN3(n7), .IN4(\ram[254][4] ), 
        .Q(n1471) );
  AOI221X1 U3266 ( .IN1(n37), .IN2(\ram[244][4] ), .IN3(n40), .IN4(
        \ram[243][4] ), .IN5(n1472), .QN(n1465) );
  AO22X1 U3267 ( .IN1(n28), .IN2(\ram[247][4] ), .IN3(n25), .IN4(\ram[248][4] ), .Q(n1472) );
  NAND4X0 U3268 ( .IN1(n1473), .IN2(n1474), .IN3(n1475), .IN4(n1476), .QN(
        n1445) );
  AOI221X1 U3269 ( .IN1(n157), .IN2(\ram[204][4] ), .IN3(n160), .IN4(
        \ram[203][4] ), .IN5(n1477), .QN(n1476) );
  AO22X1 U3270 ( .IN1(n148), .IN2(\ram[207][4] ), .IN3(n145), .IN4(
        \ram[208][4] ), .Q(n1477) );
  AOI221X1 U3271 ( .IN1(n181), .IN2(\ram[196][4] ), .IN3(n184), .IN4(
        \ram[195][4] ), .IN5(n1478), .QN(n1475) );
  AO22X1 U3272 ( .IN1(n172), .IN2(\ram[199][4] ), .IN3(n169), .IN4(
        \ram[200][4] ), .Q(n1478) );
  AOI221X1 U3273 ( .IN1(n109), .IN2(\ram[220][4] ), .IN3(n112), .IN4(
        \ram[219][4] ), .IN5(n1479), .QN(n1474) );
  AO22X1 U3274 ( .IN1(n100), .IN2(\ram[223][4] ), .IN3(n97), .IN4(
        \ram[224][4] ), .Q(n1479) );
  AOI221X1 U3275 ( .IN1(n133), .IN2(\ram[212][4] ), .IN3(n136), .IN4(
        \ram[211][4] ), .IN5(n1480), .QN(n1473) );
  AO22X1 U3276 ( .IN1(n124), .IN2(\ram[215][4] ), .IN3(n121), .IN4(
        \ram[216][4] ), .Q(n1480) );
  NAND4X0 U3278 ( .IN1(n1485), .IN2(n1486), .IN3(n1487), .IN4(n1488), .QN(
        n1484) );
  AOI221X1 U3279 ( .IN1(n637), .IN2(\ram[44][4] ), .IN3(n640), .IN4(
        \ram[43][4] ), .IN5(n1489), .QN(n1488) );
  AO22X1 U3280 ( .IN1(n628), .IN2(\ram[47][4] ), .IN3(n625), .IN4(\ram[48][4] ), .Q(n1489) );
  AOI221X1 U3281 ( .IN1(n661), .IN2(\ram[36][4] ), .IN3(n664), .IN4(
        \ram[35][4] ), .IN5(n1490), .QN(n1487) );
  AO22X1 U3282 ( .IN1(n652), .IN2(\ram[39][4] ), .IN3(n649), .IN4(\ram[40][4] ), .Q(n1490) );
  AOI221X1 U3283 ( .IN1(n589), .IN2(\ram[60][4] ), .IN3(n592), .IN4(
        \ram[59][4] ), .IN5(n1491), .QN(n1486) );
  AO22X1 U3284 ( .IN1(n580), .IN2(\ram[63][4] ), .IN3(n577), .IN4(\ram[64][4] ), .Q(n1491) );
  AOI221X1 U3285 ( .IN1(n613), .IN2(\ram[52][4] ), .IN3(n616), .IN4(
        \ram[51][4] ), .IN5(n1492), .QN(n1485) );
  AO22X1 U3286 ( .IN1(n604), .IN2(\ram[55][4] ), .IN3(n601), .IN4(\ram[56][4] ), .Q(n1492) );
  NAND4X0 U3287 ( .IN1(n1493), .IN2(n1494), .IN3(n1495), .IN4(n1496), .QN(
        n1483) );
  AOI221X1 U3288 ( .IN1(n733), .IN2(\ram[12][4] ), .IN3(n736), .IN4(
        \ram[11][4] ), .IN5(n1497), .QN(n1496) );
  AO22X1 U3289 ( .IN1(n724), .IN2(\ram[15][4] ), .IN3(n721), .IN4(\ram[16][4] ), .Q(n1497) );
  AOI221X1 U3290 ( .IN1(n757), .IN2(\ram[4][4] ), .IN3(n760), .IN4(\ram[3][4] ), .IN5(n1498), .QN(n1495) );
  AO22X1 U3291 ( .IN1(n748), .IN2(\ram[7][4] ), .IN3(n745), .IN4(\ram[8][4] ), 
        .Q(n1498) );
  AOI221X1 U3292 ( .IN1(n685), .IN2(\ram[28][4] ), .IN3(n688), .IN4(
        \ram[27][4] ), .IN5(n1499), .QN(n1494) );
  AO22X1 U3293 ( .IN1(n676), .IN2(\ram[31][4] ), .IN3(n673), .IN4(\ram[32][4] ), .Q(n1499) );
  AOI221X1 U3294 ( .IN1(n709), .IN2(\ram[20][4] ), .IN3(n712), .IN4(
        \ram[19][4] ), .IN5(n1500), .QN(n1493) );
  AO22X1 U3295 ( .IN1(n700), .IN2(\ram[23][4] ), .IN3(n697), .IN4(\ram[24][4] ), .Q(n1500) );
  NAND4X0 U3296 ( .IN1(n1501), .IN2(n1502), .IN3(n1503), .IN4(n1504), .QN(
        n1482) );
  AOI221X1 U3297 ( .IN1(n445), .IN2(\ram[108][4] ), .IN3(n448), .IN4(
        \ram[107][4] ), .IN5(n1505), .QN(n1504) );
  AO22X1 U3298 ( .IN1(n436), .IN2(\ram[111][4] ), .IN3(n433), .IN4(
        \ram[112][4] ), .Q(n1505) );
  AOI221X1 U3299 ( .IN1(n469), .IN2(\ram[100][4] ), .IN3(n472), .IN4(
        \ram[99][4] ), .IN5(n1506), .QN(n1503) );
  AO22X1 U3300 ( .IN1(n460), .IN2(\ram[103][4] ), .IN3(n457), .IN4(
        \ram[104][4] ), .Q(n1506) );
  AOI221X1 U3301 ( .IN1(n397), .IN2(\ram[124][4] ), .IN3(n400), .IN4(
        \ram[123][4] ), .IN5(n1507), .QN(n1502) );
  AO22X1 U3302 ( .IN1(n388), .IN2(\ram[127][4] ), .IN3(n385), .IN4(
        \ram[128][4] ), .Q(n1507) );
  AOI221X1 U3303 ( .IN1(n421), .IN2(\ram[116][4] ), .IN3(n424), .IN4(
        \ram[115][4] ), .IN5(n1508), .QN(n1501) );
  AO22X1 U3304 ( .IN1(n412), .IN2(\ram[119][4] ), .IN3(n409), .IN4(
        \ram[120][4] ), .Q(n1508) );
  NAND4X0 U3305 ( .IN1(n1509), .IN2(n1510), .IN3(n1511), .IN4(n1512), .QN(
        n1481) );
  AOI221X1 U3306 ( .IN1(n541), .IN2(\ram[76][4] ), .IN3(n544), .IN4(
        \ram[75][4] ), .IN5(n1513), .QN(n1512) );
  AO22X1 U3307 ( .IN1(n532), .IN2(\ram[79][4] ), .IN3(n529), .IN4(\ram[80][4] ), .Q(n1513) );
  AOI221X1 U3308 ( .IN1(n565), .IN2(\ram[68][4] ), .IN3(n568), .IN4(
        \ram[67][4] ), .IN5(n1514), .QN(n1511) );
  AO22X1 U3309 ( .IN1(n556), .IN2(\ram[71][4] ), .IN3(n553), .IN4(\ram[72][4] ), .Q(n1514) );
  AOI221X1 U3310 ( .IN1(n493), .IN2(\ram[92][4] ), .IN3(n496), .IN4(
        \ram[91][4] ), .IN5(n1515), .QN(n1510) );
  AO22X1 U3311 ( .IN1(n484), .IN2(\ram[95][4] ), .IN3(n481), .IN4(\ram[96][4] ), .Q(n1515) );
  AOI221X1 U3312 ( .IN1(n517), .IN2(\ram[84][4] ), .IN3(n520), .IN4(
        \ram[83][4] ), .IN5(n1516), .QN(n1509) );
  AO22X1 U3313 ( .IN1(n508), .IN2(\ram[87][4] ), .IN3(n505), .IN4(\ram[88][4] ), .Q(n1516) );
  AO22X1 U3314 ( .IN1(n771), .IN2(dataout[5]), .IN3(n4174), .IN4(n1517), .Q(
        n2025) );
  NAND4X0 U3315 ( .IN1(n1518), .IN2(n1519), .IN3(n1520), .IN4(n1521), .QN(
        n1517) );
  NAND4X0 U3317 ( .IN1(n1526), .IN2(n1527), .IN3(n1528), .IN4(n1529), .QN(
        n1525) );
  AOI221X1 U3318 ( .IN1(n259), .IN2(\ram[170][5] ), .IN3(n262), .IN4(
        \ram[169][5] ), .IN5(n1530), .QN(n1529) );
  AO22X1 U3319 ( .IN1(n250), .IN2(\ram[173][5] ), .IN3(n247), .IN4(
        \ram[174][5] ), .Q(n1530) );
  AOI221X1 U3320 ( .IN1(n283), .IN2(\ram[162][5] ), .IN3(n286), .IN4(
        \ram[161][5] ), .IN5(n1531), .QN(n1528) );
  AO22X1 U3321 ( .IN1(n274), .IN2(\ram[165][5] ), .IN3(n271), .IN4(
        \ram[166][5] ), .Q(n1531) );
  AOI221X1 U3322 ( .IN1(n211), .IN2(\ram[186][5] ), .IN3(n214), .IN4(
        \ram[185][5] ), .IN5(n1532), .QN(n1527) );
  AO22X1 U3323 ( .IN1(n196), .IN2(\ram[191][5] ), .IN3(n193), .IN4(
        \ram[192][5] ), .Q(n1532) );
  AOI221X1 U3324 ( .IN1(n235), .IN2(\ram[178][5] ), .IN3(n238), .IN4(
        \ram[177][5] ), .IN5(n1533), .QN(n1526) );
  AO22X1 U3325 ( .IN1(n226), .IN2(\ram[181][5] ), .IN3(n223), .IN4(
        \ram[182][5] ), .Q(n1533) );
  NAND4X0 U3326 ( .IN1(n1534), .IN2(n1535), .IN3(n1536), .IN4(n1537), .QN(
        n1524) );
  AOI221X1 U3327 ( .IN1(n355), .IN2(\ram[138][5] ), .IN3(n358), .IN4(
        \ram[137][5] ), .IN5(n1538), .QN(n1537) );
  AO22X1 U3328 ( .IN1(n346), .IN2(\ram[141][5] ), .IN3(n343), .IN4(
        \ram[142][5] ), .Q(n1538) );
  AOI221X1 U3329 ( .IN1(n379), .IN2(\ram[130][5] ), .IN3(n382), .IN4(
        \ram[129][5] ), .IN5(n1539), .QN(n1536) );
  AO22X1 U3330 ( .IN1(n370), .IN2(\ram[133][5] ), .IN3(n367), .IN4(
        \ram[134][5] ), .Q(n1539) );
  AOI221X1 U3331 ( .IN1(n307), .IN2(\ram[154][5] ), .IN3(n310), .IN4(
        \ram[153][5] ), .IN5(n1540), .QN(n1535) );
  AO22X1 U3332 ( .IN1(n298), .IN2(\ram[157][5] ), .IN3(n295), .IN4(
        \ram[158][5] ), .Q(n1540) );
  AOI221X1 U3333 ( .IN1(n331), .IN2(\ram[146][5] ), .IN3(n334), .IN4(
        \ram[145][5] ), .IN5(n1541), .QN(n1534) );
  AO22X1 U3334 ( .IN1(n322), .IN2(\ram[149][5] ), .IN3(n319), .IN4(
        \ram[150][5] ), .Q(n1541) );
  NAND4X0 U3335 ( .IN1(n1542), .IN2(n1543), .IN3(n1544), .IN4(n1545), .QN(
        n1523) );
  AOI221X1 U3336 ( .IN1(n70), .IN2(\ram[233][5] ), .IN3(n49), .IN4(
        \ram[240][5] ), .IN5(n1546), .QN(n1545) );
  AO22X1 U3337 ( .IN1(n139), .IN2(\ram[210][5] ), .IN3(n52), .IN4(
        \ram[239][5] ), .Q(n1546) );
  AOI221X1 U3338 ( .IN1(n94), .IN2(\ram[225][5] ), .IN3(n79), .IN4(
        \ram[230][5] ), .IN5(n1547), .QN(n1544) );
  AO22X1 U3339 ( .IN1(n67), .IN2(\ram[234][5] ), .IN3(n82), .IN4(\ram[229][5] ), .Q(n1547) );
  AOI221X1 U3340 ( .IN1(n13), .IN2(\ram[252][5] ), .IN3(n16), .IN4(
        \ram[251][5] ), .IN5(n1548), .QN(n1543) );
  AO22X1 U3341 ( .IN1(n91), .IN2(\ram[226][5] ), .IN3(n3), .IN4(\ram[255][5] ), 
        .Q(n1548) );
  AOI221X1 U3342 ( .IN1(n43), .IN2(\ram[242][5] ), .IN3(n46), .IN4(
        \ram[241][5] ), .IN5(n1549), .QN(n1542) );
  AO22X1 U3343 ( .IN1(n34), .IN2(\ram[245][5] ), .IN3(n31), .IN4(\ram[246][5] ), .Q(n1549) );
  NAND4X0 U3344 ( .IN1(n1550), .IN2(n1551), .IN3(n1552), .IN4(n1553), .QN(
        n1522) );
  AOI221X1 U3345 ( .IN1(n166), .IN2(\ram[201][5] ), .IN3(n151), .IN4(
        \ram[206][5] ), .IN5(n1554), .QN(n1553) );
  AO22X1 U3346 ( .IN1(n769), .IN2(\ram[0][5] ), .IN3(n154), .IN4(\ram[205][5] ), .Q(n1554) );
  AOI221X1 U3347 ( .IN1(n190), .IN2(\ram[193][5] ), .IN3(n175), .IN4(
        \ram[198][5] ), .IN5(n1555), .QN(n1552) );
  AO22X1 U3348 ( .IN1(n163), .IN2(\ram[202][5] ), .IN3(n178), .IN4(
        \ram[197][5] ), .Q(n1555) );
  AOI221X1 U3349 ( .IN1(n106), .IN2(\ram[221][5] ), .IN3(n187), .IN4(
        \ram[194][5] ), .IN5(n1556), .QN(n1551) );
  AO22X1 U3350 ( .IN1(n103), .IN2(\ram[222][5] ), .IN3(n118), .IN4(
        \ram[217][5] ), .Q(n1556) );
  AOI221X1 U3351 ( .IN1(n142), .IN2(\ram[209][5] ), .IN3(n127), .IN4(
        \ram[214][5] ), .IN5(n1557), .QN(n1550) );
  AO22X1 U3352 ( .IN1(n115), .IN2(\ram[218][5] ), .IN3(n130), .IN4(
        \ram[213][5] ), .Q(n1557) );
  NAND4X0 U3354 ( .IN1(n1562), .IN2(n1563), .IN3(n1564), .IN4(n1565), .QN(
        n1561) );
  AOI221X1 U3355 ( .IN1(n643), .IN2(\ram[42][5] ), .IN3(n646), .IN4(
        \ram[41][5] ), .IN5(n1566), .QN(n1565) );
  AO22X1 U3356 ( .IN1(n634), .IN2(\ram[45][5] ), .IN3(n631), .IN4(\ram[46][5] ), .Q(n1566) );
  AOI221X1 U3357 ( .IN1(n667), .IN2(\ram[34][5] ), .IN3(n670), .IN4(
        \ram[33][5] ), .IN5(n1567), .QN(n1564) );
  AO22X1 U3358 ( .IN1(n658), .IN2(\ram[37][5] ), .IN3(n655), .IN4(\ram[38][5] ), .Q(n1567) );
  AOI221X1 U3359 ( .IN1(n595), .IN2(\ram[58][5] ), .IN3(n598), .IN4(
        \ram[57][5] ), .IN5(n1568), .QN(n1563) );
  AO22X1 U3360 ( .IN1(n586), .IN2(\ram[61][5] ), .IN3(n583), .IN4(\ram[62][5] ), .Q(n1568) );
  AOI221X1 U3361 ( .IN1(n619), .IN2(\ram[50][5] ), .IN3(n622), .IN4(
        \ram[49][5] ), .IN5(n1569), .QN(n1562) );
  AO22X1 U3362 ( .IN1(n610), .IN2(\ram[53][5] ), .IN3(n607), .IN4(\ram[54][5] ), .Q(n1569) );
  NAND4X0 U3363 ( .IN1(n1570), .IN2(n1571), .IN3(n1572), .IN4(n1573), .QN(
        n1560) );
  AOI221X1 U3364 ( .IN1(n739), .IN2(\ram[10][5] ), .IN3(n742), .IN4(
        \ram[9][5] ), .IN5(n1574), .QN(n1573) );
  AO22X1 U3365 ( .IN1(n730), .IN2(\ram[13][5] ), .IN3(n727), .IN4(\ram[14][5] ), .Q(n1574) );
  AOI221X1 U3366 ( .IN1(n763), .IN2(\ram[2][5] ), .IN3(n766), .IN4(\ram[1][5] ), .IN5(n1575), .QN(n1572) );
  AO22X1 U3367 ( .IN1(n754), .IN2(\ram[5][5] ), .IN3(n751), .IN4(\ram[6][5] ), 
        .Q(n1575) );
  AOI221X1 U3368 ( .IN1(n691), .IN2(\ram[26][5] ), .IN3(n694), .IN4(
        \ram[25][5] ), .IN5(n1576), .QN(n1571) );
  AO22X1 U3369 ( .IN1(n682), .IN2(\ram[29][5] ), .IN3(n679), .IN4(\ram[30][5] ), .Q(n1576) );
  AOI221X1 U3370 ( .IN1(n715), .IN2(\ram[18][5] ), .IN3(n718), .IN4(
        \ram[17][5] ), .IN5(n1577), .QN(n1570) );
  AO22X1 U3371 ( .IN1(n706), .IN2(\ram[21][5] ), .IN3(n703), .IN4(\ram[22][5] ), .Q(n1577) );
  NAND4X0 U3372 ( .IN1(n1578), .IN2(n1579), .IN3(n1580), .IN4(n1581), .QN(
        n1559) );
  AOI221X1 U3373 ( .IN1(n451), .IN2(\ram[106][5] ), .IN3(n454), .IN4(
        \ram[105][5] ), .IN5(n1582), .QN(n1581) );
  AO22X1 U3374 ( .IN1(n442), .IN2(\ram[109][5] ), .IN3(n439), .IN4(
        \ram[110][5] ), .Q(n1582) );
  AOI221X1 U3375 ( .IN1(n475), .IN2(\ram[98][5] ), .IN3(n478), .IN4(
        \ram[97][5] ), .IN5(n1583), .QN(n1580) );
  AO22X1 U3376 ( .IN1(n466), .IN2(\ram[101][5] ), .IN3(n463), .IN4(
        \ram[102][5] ), .Q(n1583) );
  AOI221X1 U3377 ( .IN1(n403), .IN2(\ram[122][5] ), .IN3(n406), .IN4(
        \ram[121][5] ), .IN5(n1584), .QN(n1579) );
  AO22X1 U3378 ( .IN1(n394), .IN2(\ram[125][5] ), .IN3(n391), .IN4(
        \ram[126][5] ), .Q(n1584) );
  AOI221X1 U3379 ( .IN1(n427), .IN2(\ram[114][5] ), .IN3(n430), .IN4(
        \ram[113][5] ), .IN5(n1585), .QN(n1578) );
  AO22X1 U3380 ( .IN1(n418), .IN2(\ram[117][5] ), .IN3(n415), .IN4(
        \ram[118][5] ), .Q(n1585) );
  NAND4X0 U3381 ( .IN1(n1586), .IN2(n1587), .IN3(n1588), .IN4(n1589), .QN(
        n1558) );
  AOI221X1 U3382 ( .IN1(n547), .IN2(\ram[74][5] ), .IN3(n550), .IN4(
        \ram[73][5] ), .IN5(n1590), .QN(n1589) );
  AO22X1 U3383 ( .IN1(n538), .IN2(\ram[77][5] ), .IN3(n535), .IN4(\ram[78][5] ), .Q(n1590) );
  AOI221X1 U3384 ( .IN1(n571), .IN2(\ram[66][5] ), .IN3(n574), .IN4(
        \ram[65][5] ), .IN5(n1591), .QN(n1588) );
  AO22X1 U3385 ( .IN1(n562), .IN2(\ram[69][5] ), .IN3(n559), .IN4(\ram[70][5] ), .Q(n1591) );
  AOI221X1 U3386 ( .IN1(n499), .IN2(\ram[90][5] ), .IN3(n502), .IN4(
        \ram[89][5] ), .IN5(n1592), .QN(n1587) );
  AO22X1 U3387 ( .IN1(n490), .IN2(\ram[93][5] ), .IN3(n487), .IN4(\ram[94][5] ), .Q(n1592) );
  AOI221X1 U3388 ( .IN1(n523), .IN2(\ram[82][5] ), .IN3(n526), .IN4(
        \ram[81][5] ), .IN5(n1593), .QN(n1586) );
  AO22X1 U3389 ( .IN1(n514), .IN2(\ram[85][5] ), .IN3(n511), .IN4(\ram[86][5] ), .Q(n1593) );
  NAND4X0 U3391 ( .IN1(n1598), .IN2(n1599), .IN3(n1600), .IN4(n1601), .QN(
        n1597) );
  AOI221X1 U3392 ( .IN1(n253), .IN2(\ram[172][5] ), .IN3(n256), .IN4(
        \ram[171][5] ), .IN5(n1602), .QN(n1601) );
  AO22X1 U3393 ( .IN1(n244), .IN2(\ram[175][5] ), .IN3(n241), .IN4(
        \ram[176][5] ), .Q(n1602) );
  AOI221X1 U3394 ( .IN1(n277), .IN2(\ram[164][5] ), .IN3(n280), .IN4(
        \ram[163][5] ), .IN5(n1603), .QN(n1600) );
  AO22X1 U3395 ( .IN1(n268), .IN2(\ram[167][5] ), .IN3(n265), .IN4(
        \ram[168][5] ), .Q(n1603) );
  AOI221X1 U3396 ( .IN1(n205), .IN2(\ram[188][5] ), .IN3(n208), .IN4(
        \ram[187][5] ), .IN5(n1604), .QN(n1599) );
  AO22X1 U3397 ( .IN1(n202), .IN2(\ram[189][5] ), .IN3(n199), .IN4(
        \ram[190][5] ), .Q(n1604) );
  AOI221X1 U3398 ( .IN1(n229), .IN2(\ram[180][5] ), .IN3(n232), .IN4(
        \ram[179][5] ), .IN5(n1605), .QN(n1598) );
  AO22X1 U3399 ( .IN1(n220), .IN2(\ram[183][5] ), .IN3(n217), .IN4(
        \ram[184][5] ), .Q(n1605) );
  NAND4X0 U3400 ( .IN1(n1606), .IN2(n1607), .IN3(n1608), .IN4(n1609), .QN(
        n1596) );
  AOI221X1 U3401 ( .IN1(n349), .IN2(\ram[140][5] ), .IN3(n352), .IN4(
        \ram[139][5] ), .IN5(n1610), .QN(n1609) );
  AO22X1 U3402 ( .IN1(n340), .IN2(\ram[143][5] ), .IN3(n337), .IN4(
        \ram[144][5] ), .Q(n1610) );
  AOI221X1 U3403 ( .IN1(n373), .IN2(\ram[132][5] ), .IN3(n376), .IN4(
        \ram[131][5] ), .IN5(n1611), .QN(n1608) );
  AO22X1 U3404 ( .IN1(n364), .IN2(\ram[135][5] ), .IN3(n361), .IN4(
        \ram[136][5] ), .Q(n1611) );
  AOI221X1 U3405 ( .IN1(n301), .IN2(\ram[156][5] ), .IN3(n304), .IN4(
        \ram[155][5] ), .IN5(n1612), .QN(n1607) );
  AO22X1 U3406 ( .IN1(n292), .IN2(\ram[159][5] ), .IN3(n289), .IN4(
        \ram[160][5] ), .Q(n1612) );
  AOI221X1 U3407 ( .IN1(n325), .IN2(\ram[148][5] ), .IN3(n328), .IN4(
        \ram[147][5] ), .IN5(n1613), .QN(n1606) );
  AO22X1 U3408 ( .IN1(n316), .IN2(\ram[151][5] ), .IN3(n313), .IN4(
        \ram[152][5] ), .Q(n1613) );
  NAND4X0 U3409 ( .IN1(n1614), .IN2(n1615), .IN3(n1616), .IN4(n1617), .QN(
        n1595) );
  AOI221X1 U3410 ( .IN1(n61), .IN2(\ram[236][5] ), .IN3(n64), .IN4(
        \ram[235][5] ), .IN5(n1618), .QN(n1617) );
  AO22X1 U3411 ( .IN1(n58), .IN2(\ram[237][5] ), .IN3(n55), .IN4(\ram[238][5] ), .Q(n1618) );
  AOI221X1 U3412 ( .IN1(n85), .IN2(\ram[228][5] ), .IN3(n88), .IN4(
        \ram[227][5] ), .IN5(n1619), .QN(n1616) );
  AO22X1 U3413 ( .IN1(n76), .IN2(\ram[231][5] ), .IN3(n73), .IN4(\ram[232][5] ), .Q(n1619) );
  AOI221X1 U3414 ( .IN1(n19), .IN2(\ram[250][5] ), .IN3(n22), .IN4(
        \ram[249][5] ), .IN5(n1620), .QN(n1615) );
  AO22X1 U3415 ( .IN1(n10), .IN2(\ram[253][5] ), .IN3(n7), .IN4(\ram[254][5] ), 
        .Q(n1620) );
  AOI221X1 U3416 ( .IN1(n37), .IN2(\ram[244][5] ), .IN3(n40), .IN4(
        \ram[243][5] ), .IN5(n1621), .QN(n1614) );
  AO22X1 U3417 ( .IN1(n28), .IN2(\ram[247][5] ), .IN3(n25), .IN4(\ram[248][5] ), .Q(n1621) );
  NAND4X0 U3418 ( .IN1(n1622), .IN2(n1623), .IN3(n1624), .IN4(n1625), .QN(
        n1594) );
  AOI221X1 U3419 ( .IN1(n157), .IN2(\ram[204][5] ), .IN3(n160), .IN4(
        \ram[203][5] ), .IN5(n1626), .QN(n1625) );
  AO22X1 U3420 ( .IN1(n148), .IN2(\ram[207][5] ), .IN3(n145), .IN4(
        \ram[208][5] ), .Q(n1626) );
  AOI221X1 U3421 ( .IN1(n181), .IN2(\ram[196][5] ), .IN3(n184), .IN4(
        \ram[195][5] ), .IN5(n1627), .QN(n1624) );
  AO22X1 U3422 ( .IN1(n172), .IN2(\ram[199][5] ), .IN3(n169), .IN4(
        \ram[200][5] ), .Q(n1627) );
  AOI221X1 U3423 ( .IN1(n109), .IN2(\ram[220][5] ), .IN3(n112), .IN4(
        \ram[219][5] ), .IN5(n1628), .QN(n1623) );
  AO22X1 U3424 ( .IN1(n100), .IN2(\ram[223][5] ), .IN3(n97), .IN4(
        \ram[224][5] ), .Q(n1628) );
  AOI221X1 U3425 ( .IN1(n133), .IN2(\ram[212][5] ), .IN3(n136), .IN4(
        \ram[211][5] ), .IN5(n1629), .QN(n1622) );
  AO22X1 U3426 ( .IN1(n124), .IN2(\ram[215][5] ), .IN3(n121), .IN4(
        \ram[216][5] ), .Q(n1629) );
  NAND4X0 U3428 ( .IN1(n1634), .IN2(n1635), .IN3(n1636), .IN4(n1637), .QN(
        n1633) );
  AOI221X1 U3429 ( .IN1(n637), .IN2(\ram[44][5] ), .IN3(n640), .IN4(
        \ram[43][5] ), .IN5(n1638), .QN(n1637) );
  AO22X1 U3430 ( .IN1(n628), .IN2(\ram[47][5] ), .IN3(n625), .IN4(\ram[48][5] ), .Q(n1638) );
  AOI221X1 U3431 ( .IN1(n661), .IN2(\ram[36][5] ), .IN3(n664), .IN4(
        \ram[35][5] ), .IN5(n1639), .QN(n1636) );
  AO22X1 U3432 ( .IN1(n652), .IN2(\ram[39][5] ), .IN3(n649), .IN4(\ram[40][5] ), .Q(n1639) );
  AOI221X1 U3433 ( .IN1(n589), .IN2(\ram[60][5] ), .IN3(n592), .IN4(
        \ram[59][5] ), .IN5(n1640), .QN(n1635) );
  AO22X1 U3434 ( .IN1(n580), .IN2(\ram[63][5] ), .IN3(n577), .IN4(\ram[64][5] ), .Q(n1640) );
  AOI221X1 U3435 ( .IN1(n613), .IN2(\ram[52][5] ), .IN3(n616), .IN4(
        \ram[51][5] ), .IN5(n1641), .QN(n1634) );
  AO22X1 U3436 ( .IN1(n604), .IN2(\ram[55][5] ), .IN3(n601), .IN4(\ram[56][5] ), .Q(n1641) );
  NAND4X0 U3437 ( .IN1(n1642), .IN2(n1643), .IN3(n1644), .IN4(n1645), .QN(
        n1632) );
  AOI221X1 U3438 ( .IN1(n733), .IN2(\ram[12][5] ), .IN3(n736), .IN4(
        \ram[11][5] ), .IN5(n1646), .QN(n1645) );
  AO22X1 U3439 ( .IN1(n724), .IN2(\ram[15][5] ), .IN3(n721), .IN4(\ram[16][5] ), .Q(n1646) );
  AOI221X1 U3440 ( .IN1(n757), .IN2(\ram[4][5] ), .IN3(n760), .IN4(\ram[3][5] ), .IN5(n1647), .QN(n1644) );
  AO22X1 U3441 ( .IN1(n748), .IN2(\ram[7][5] ), .IN3(n745), .IN4(\ram[8][5] ), 
        .Q(n1647) );
  AOI221X1 U3442 ( .IN1(n685), .IN2(\ram[28][5] ), .IN3(n688), .IN4(
        \ram[27][5] ), .IN5(n1648), .QN(n1643) );
  AO22X1 U3443 ( .IN1(n676), .IN2(\ram[31][5] ), .IN3(n673), .IN4(\ram[32][5] ), .Q(n1648) );
  AOI221X1 U3444 ( .IN1(n709), .IN2(\ram[20][5] ), .IN3(n712), .IN4(
        \ram[19][5] ), .IN5(n1649), .QN(n1642) );
  AO22X1 U3445 ( .IN1(n700), .IN2(\ram[23][5] ), .IN3(n697), .IN4(\ram[24][5] ), .Q(n1649) );
  NAND4X0 U3446 ( .IN1(n1650), .IN2(n1651), .IN3(n1652), .IN4(n1653), .QN(
        n1631) );
  AOI221X1 U3447 ( .IN1(n445), .IN2(\ram[108][5] ), .IN3(n448), .IN4(
        \ram[107][5] ), .IN5(n1654), .QN(n1653) );
  AO22X1 U3448 ( .IN1(n436), .IN2(\ram[111][5] ), .IN3(n433), .IN4(
        \ram[112][5] ), .Q(n1654) );
  AOI221X1 U3449 ( .IN1(n469), .IN2(\ram[100][5] ), .IN3(n472), .IN4(
        \ram[99][5] ), .IN5(n1655), .QN(n1652) );
  AO22X1 U3450 ( .IN1(n460), .IN2(\ram[103][5] ), .IN3(n457), .IN4(
        \ram[104][5] ), .Q(n1655) );
  AOI221X1 U3451 ( .IN1(n397), .IN2(\ram[124][5] ), .IN3(n400), .IN4(
        \ram[123][5] ), .IN5(n1656), .QN(n1651) );
  AO22X1 U3452 ( .IN1(n388), .IN2(\ram[127][5] ), .IN3(n385), .IN4(
        \ram[128][5] ), .Q(n1656) );
  AOI221X1 U3453 ( .IN1(n421), .IN2(\ram[116][5] ), .IN3(n424), .IN4(
        \ram[115][5] ), .IN5(n1657), .QN(n1650) );
  AO22X1 U3454 ( .IN1(n412), .IN2(\ram[119][5] ), .IN3(n409), .IN4(
        \ram[120][5] ), .Q(n1657) );
  NAND4X0 U3455 ( .IN1(n1658), .IN2(n1659), .IN3(n1660), .IN4(n1661), .QN(
        n1630) );
  AOI221X1 U3456 ( .IN1(n541), .IN2(\ram[76][5] ), .IN3(n544), .IN4(
        \ram[75][5] ), .IN5(n1662), .QN(n1661) );
  AO22X1 U3457 ( .IN1(n532), .IN2(\ram[79][5] ), .IN3(n529), .IN4(\ram[80][5] ), .Q(n1662) );
  AOI221X1 U3458 ( .IN1(n565), .IN2(\ram[68][5] ), .IN3(n568), .IN4(
        \ram[67][5] ), .IN5(n1663), .QN(n1660) );
  AO22X1 U3459 ( .IN1(n556), .IN2(\ram[71][5] ), .IN3(n553), .IN4(\ram[72][5] ), .Q(n1663) );
  AOI221X1 U3460 ( .IN1(n493), .IN2(\ram[92][5] ), .IN3(n496), .IN4(
        \ram[91][5] ), .IN5(n1664), .QN(n1659) );
  AO22X1 U3461 ( .IN1(n484), .IN2(\ram[95][5] ), .IN3(n481), .IN4(\ram[96][5] ), .Q(n1664) );
  AOI221X1 U3462 ( .IN1(n517), .IN2(\ram[84][5] ), .IN3(n520), .IN4(
        \ram[83][5] ), .IN5(n1665), .QN(n1658) );
  AO22X1 U3463 ( .IN1(n508), .IN2(\ram[87][5] ), .IN3(n505), .IN4(\ram[88][5] ), .Q(n1665) );
  AO22X1 U3464 ( .IN1(n771), .IN2(dataout[6]), .IN3(n4174), .IN4(n1666), .Q(
        n2026) );
  NAND4X0 U3465 ( .IN1(n1667), .IN2(n1668), .IN3(n1669), .IN4(n1670), .QN(
        n1666) );
  NAND4X0 U3467 ( .IN1(n1675), .IN2(n1676), .IN3(n1677), .IN4(n1678), .QN(
        n1674) );
  AOI221X1 U3468 ( .IN1(n259), .IN2(\ram[170][6] ), .IN3(n262), .IN4(
        \ram[169][6] ), .IN5(n1679), .QN(n1678) );
  AO22X1 U3469 ( .IN1(n250), .IN2(\ram[173][6] ), .IN3(n247), .IN4(
        \ram[174][6] ), .Q(n1679) );
  AOI221X1 U3470 ( .IN1(n283), .IN2(\ram[162][6] ), .IN3(n286), .IN4(
        \ram[161][6] ), .IN5(n1680), .QN(n1677) );
  AO22X1 U3471 ( .IN1(n274), .IN2(\ram[165][6] ), .IN3(n271), .IN4(
        \ram[166][6] ), .Q(n1680) );
  AOI221X1 U3472 ( .IN1(n211), .IN2(\ram[186][6] ), .IN3(n214), .IN4(
        \ram[185][6] ), .IN5(n1681), .QN(n1676) );
  AO22X1 U3473 ( .IN1(n196), .IN2(\ram[191][6] ), .IN3(n193), .IN4(
        \ram[192][6] ), .Q(n1681) );
  AOI221X1 U3474 ( .IN1(n235), .IN2(\ram[178][6] ), .IN3(n238), .IN4(
        \ram[177][6] ), .IN5(n1682), .QN(n1675) );
  AO22X1 U3475 ( .IN1(n226), .IN2(\ram[181][6] ), .IN3(n223), .IN4(
        \ram[182][6] ), .Q(n1682) );
  NAND4X0 U3476 ( .IN1(n1683), .IN2(n1684), .IN3(n1685), .IN4(n1686), .QN(
        n1673) );
  AOI221X1 U3477 ( .IN1(n355), .IN2(\ram[138][6] ), .IN3(n358), .IN4(
        \ram[137][6] ), .IN5(n1687), .QN(n1686) );
  AO22X1 U3478 ( .IN1(n346), .IN2(\ram[141][6] ), .IN3(n343), .IN4(
        \ram[142][6] ), .Q(n1687) );
  AOI221X1 U3479 ( .IN1(n379), .IN2(\ram[130][6] ), .IN3(n382), .IN4(
        \ram[129][6] ), .IN5(n1688), .QN(n1685) );
  AO22X1 U3480 ( .IN1(n370), .IN2(\ram[133][6] ), .IN3(n367), .IN4(
        \ram[134][6] ), .Q(n1688) );
  AOI221X1 U3481 ( .IN1(n307), .IN2(\ram[154][6] ), .IN3(n310), .IN4(
        \ram[153][6] ), .IN5(n1689), .QN(n1684) );
  AO22X1 U3482 ( .IN1(n298), .IN2(\ram[157][6] ), .IN3(n295), .IN4(
        \ram[158][6] ), .Q(n1689) );
  AOI221X1 U3483 ( .IN1(n331), .IN2(\ram[146][6] ), .IN3(n334), .IN4(
        \ram[145][6] ), .IN5(n1690), .QN(n1683) );
  AO22X1 U3484 ( .IN1(n322), .IN2(\ram[149][6] ), .IN3(n319), .IN4(
        \ram[150][6] ), .Q(n1690) );
  NAND4X0 U3485 ( .IN1(n1691), .IN2(n1692), .IN3(n1693), .IN4(n1694), .QN(
        n1672) );
  AOI221X1 U3486 ( .IN1(n70), .IN2(\ram[233][6] ), .IN3(n49), .IN4(
        \ram[240][6] ), .IN5(n1695), .QN(n1694) );
  AO22X1 U3487 ( .IN1(n139), .IN2(\ram[210][6] ), .IN3(n52), .IN4(
        \ram[239][6] ), .Q(n1695) );
  AOI221X1 U3488 ( .IN1(n94), .IN2(\ram[225][6] ), .IN3(n79), .IN4(
        \ram[230][6] ), .IN5(n1696), .QN(n1693) );
  AO22X1 U3489 ( .IN1(n67), .IN2(\ram[234][6] ), .IN3(n82), .IN4(\ram[229][6] ), .Q(n1696) );
  AOI221X1 U3490 ( .IN1(n13), .IN2(\ram[252][6] ), .IN3(n16), .IN4(
        \ram[251][6] ), .IN5(n1697), .QN(n1692) );
  AO22X1 U3491 ( .IN1(n91), .IN2(\ram[226][6] ), .IN3(n3), .IN4(\ram[255][6] ), 
        .Q(n1697) );
  AOI221X1 U3492 ( .IN1(n43), .IN2(\ram[242][6] ), .IN3(n46), .IN4(
        \ram[241][6] ), .IN5(n1698), .QN(n1691) );
  AO22X1 U3493 ( .IN1(n34), .IN2(\ram[245][6] ), .IN3(n31), .IN4(\ram[246][6] ), .Q(n1698) );
  NAND4X0 U3494 ( .IN1(n1699), .IN2(n1700), .IN3(n1701), .IN4(n1702), .QN(
        n1671) );
  AOI221X1 U3495 ( .IN1(n166), .IN2(\ram[201][6] ), .IN3(n151), .IN4(
        \ram[206][6] ), .IN5(n1703), .QN(n1702) );
  AO22X1 U3496 ( .IN1(n769), .IN2(\ram[0][6] ), .IN3(n154), .IN4(\ram[205][6] ), .Q(n1703) );
  AOI221X1 U3497 ( .IN1(n190), .IN2(\ram[193][6] ), .IN3(n175), .IN4(
        \ram[198][6] ), .IN5(n1704), .QN(n1701) );
  AO22X1 U3498 ( .IN1(n163), .IN2(\ram[202][6] ), .IN3(n178), .IN4(
        \ram[197][6] ), .Q(n1704) );
  AOI221X1 U3499 ( .IN1(n106), .IN2(\ram[221][6] ), .IN3(n187), .IN4(
        \ram[194][6] ), .IN5(n1705), .QN(n1700) );
  AO22X1 U3500 ( .IN1(n103), .IN2(\ram[222][6] ), .IN3(n118), .IN4(
        \ram[217][6] ), .Q(n1705) );
  AOI221X1 U3501 ( .IN1(n142), .IN2(\ram[209][6] ), .IN3(n127), .IN4(
        \ram[214][6] ), .IN5(n1706), .QN(n1699) );
  AO22X1 U3502 ( .IN1(n115), .IN2(\ram[218][6] ), .IN3(n130), .IN4(
        \ram[213][6] ), .Q(n1706) );
  NAND4X0 U3504 ( .IN1(n1711), .IN2(n1712), .IN3(n1713), .IN4(n1714), .QN(
        n1710) );
  AOI221X1 U3505 ( .IN1(n643), .IN2(\ram[42][6] ), .IN3(n646), .IN4(
        \ram[41][6] ), .IN5(n1715), .QN(n1714) );
  AO22X1 U3506 ( .IN1(n634), .IN2(\ram[45][6] ), .IN3(n631), .IN4(\ram[46][6] ), .Q(n1715) );
  AOI221X1 U3507 ( .IN1(n667), .IN2(\ram[34][6] ), .IN3(n670), .IN4(
        \ram[33][6] ), .IN5(n1716), .QN(n1713) );
  AO22X1 U3508 ( .IN1(n658), .IN2(\ram[37][6] ), .IN3(n655), .IN4(\ram[38][6] ), .Q(n1716) );
  AOI221X1 U3509 ( .IN1(n595), .IN2(\ram[58][6] ), .IN3(n598), .IN4(
        \ram[57][6] ), .IN5(n1717), .QN(n1712) );
  AO22X1 U3510 ( .IN1(n586), .IN2(\ram[61][6] ), .IN3(n583), .IN4(\ram[62][6] ), .Q(n1717) );
  AOI221X1 U3511 ( .IN1(n619), .IN2(\ram[50][6] ), .IN3(n622), .IN4(
        \ram[49][6] ), .IN5(n1718), .QN(n1711) );
  AO22X1 U3512 ( .IN1(n610), .IN2(\ram[53][6] ), .IN3(n607), .IN4(\ram[54][6] ), .Q(n1718) );
  NAND4X0 U3513 ( .IN1(n1719), .IN2(n1720), .IN3(n1721), .IN4(n1722), .QN(
        n1709) );
  AOI221X1 U3514 ( .IN1(n739), .IN2(\ram[10][6] ), .IN3(n742), .IN4(
        \ram[9][6] ), .IN5(n1723), .QN(n1722) );
  AO22X1 U3515 ( .IN1(n730), .IN2(\ram[13][6] ), .IN3(n727), .IN4(\ram[14][6] ), .Q(n1723) );
  AOI221X1 U3516 ( .IN1(n763), .IN2(\ram[2][6] ), .IN3(n766), .IN4(\ram[1][6] ), .IN5(n1724), .QN(n1721) );
  AO22X1 U3517 ( .IN1(n754), .IN2(\ram[5][6] ), .IN3(n751), .IN4(\ram[6][6] ), 
        .Q(n1724) );
  AOI221X1 U3518 ( .IN1(n691), .IN2(\ram[26][6] ), .IN3(n694), .IN4(
        \ram[25][6] ), .IN5(n1725), .QN(n1720) );
  AO22X1 U3519 ( .IN1(n682), .IN2(\ram[29][6] ), .IN3(n679), .IN4(\ram[30][6] ), .Q(n1725) );
  AOI221X1 U3520 ( .IN1(n715), .IN2(\ram[18][6] ), .IN3(n718), .IN4(
        \ram[17][6] ), .IN5(n1726), .QN(n1719) );
  AO22X1 U3521 ( .IN1(n706), .IN2(\ram[21][6] ), .IN3(n703), .IN4(\ram[22][6] ), .Q(n1726) );
  NAND4X0 U3522 ( .IN1(n1727), .IN2(n1728), .IN3(n1729), .IN4(n1730), .QN(
        n1708) );
  AOI221X1 U3523 ( .IN1(n451), .IN2(\ram[106][6] ), .IN3(n454), .IN4(
        \ram[105][6] ), .IN5(n1731), .QN(n1730) );
  AO22X1 U3524 ( .IN1(n442), .IN2(\ram[109][6] ), .IN3(n439), .IN4(
        \ram[110][6] ), .Q(n1731) );
  AOI221X1 U3525 ( .IN1(n475), .IN2(\ram[98][6] ), .IN3(n478), .IN4(
        \ram[97][6] ), .IN5(n1732), .QN(n1729) );
  AO22X1 U3526 ( .IN1(n466), .IN2(\ram[101][6] ), .IN3(n463), .IN4(
        \ram[102][6] ), .Q(n1732) );
  AOI221X1 U3527 ( .IN1(n403), .IN2(\ram[122][6] ), .IN3(n406), .IN4(
        \ram[121][6] ), .IN5(n1733), .QN(n1728) );
  AO22X1 U3528 ( .IN1(n394), .IN2(\ram[125][6] ), .IN3(n391), .IN4(
        \ram[126][6] ), .Q(n1733) );
  AOI221X1 U3529 ( .IN1(n427), .IN2(\ram[114][6] ), .IN3(n430), .IN4(
        \ram[113][6] ), .IN5(n1734), .QN(n1727) );
  AO22X1 U3530 ( .IN1(n418), .IN2(\ram[117][6] ), .IN3(n415), .IN4(
        \ram[118][6] ), .Q(n1734) );
  NAND4X0 U3531 ( .IN1(n1735), .IN2(n1736), .IN3(n1737), .IN4(n1738), .QN(
        n1707) );
  AOI221X1 U3532 ( .IN1(n547), .IN2(\ram[74][6] ), .IN3(n550), .IN4(
        \ram[73][6] ), .IN5(n1739), .QN(n1738) );
  AO22X1 U3533 ( .IN1(n538), .IN2(\ram[77][6] ), .IN3(n535), .IN4(\ram[78][6] ), .Q(n1739) );
  AOI221X1 U3534 ( .IN1(n571), .IN2(\ram[66][6] ), .IN3(n574), .IN4(
        \ram[65][6] ), .IN5(n1740), .QN(n1737) );
  AO22X1 U3535 ( .IN1(n562), .IN2(\ram[69][6] ), .IN3(n559), .IN4(\ram[70][6] ), .Q(n1740) );
  AOI221X1 U3536 ( .IN1(n499), .IN2(\ram[90][6] ), .IN3(n502), .IN4(
        \ram[89][6] ), .IN5(n1741), .QN(n1736) );
  AO22X1 U3537 ( .IN1(n490), .IN2(\ram[93][6] ), .IN3(n487), .IN4(\ram[94][6] ), .Q(n1741) );
  AOI221X1 U3538 ( .IN1(n523), .IN2(\ram[82][6] ), .IN3(n526), .IN4(
        \ram[81][6] ), .IN5(n1742), .QN(n1735) );
  AO22X1 U3539 ( .IN1(n514), .IN2(\ram[85][6] ), .IN3(n511), .IN4(\ram[86][6] ), .Q(n1742) );
  NAND4X0 U3541 ( .IN1(n1747), .IN2(n1748), .IN3(n1749), .IN4(n1750), .QN(
        n1746) );
  AOI221X1 U3542 ( .IN1(n253), .IN2(\ram[172][6] ), .IN3(n256), .IN4(
        \ram[171][6] ), .IN5(n1751), .QN(n1750) );
  AO22X1 U3543 ( .IN1(n244), .IN2(\ram[175][6] ), .IN3(n241), .IN4(
        \ram[176][6] ), .Q(n1751) );
  AOI221X1 U3544 ( .IN1(n277), .IN2(\ram[164][6] ), .IN3(n280), .IN4(
        \ram[163][6] ), .IN5(n1752), .QN(n1749) );
  AO22X1 U3545 ( .IN1(n268), .IN2(\ram[167][6] ), .IN3(n265), .IN4(
        \ram[168][6] ), .Q(n1752) );
  AOI221X1 U3546 ( .IN1(n205), .IN2(\ram[188][6] ), .IN3(n208), .IN4(
        \ram[187][6] ), .IN5(n1753), .QN(n1748) );
  AO22X1 U3547 ( .IN1(n202), .IN2(\ram[189][6] ), .IN3(n199), .IN4(
        \ram[190][6] ), .Q(n1753) );
  AOI221X1 U3548 ( .IN1(n229), .IN2(\ram[180][6] ), .IN3(n232), .IN4(
        \ram[179][6] ), .IN5(n1754), .QN(n1747) );
  AO22X1 U3549 ( .IN1(n220), .IN2(\ram[183][6] ), .IN3(n217), .IN4(
        \ram[184][6] ), .Q(n1754) );
  NAND4X0 U3550 ( .IN1(n1755), .IN2(n1756), .IN3(n1757), .IN4(n1758), .QN(
        n1745) );
  AOI221X1 U3551 ( .IN1(n349), .IN2(\ram[140][6] ), .IN3(n352), .IN4(
        \ram[139][6] ), .IN5(n1759), .QN(n1758) );
  AO22X1 U3552 ( .IN1(n340), .IN2(\ram[143][6] ), .IN3(n337), .IN4(
        \ram[144][6] ), .Q(n1759) );
  AOI221X1 U3553 ( .IN1(n373), .IN2(\ram[132][6] ), .IN3(n376), .IN4(
        \ram[131][6] ), .IN5(n1760), .QN(n1757) );
  AO22X1 U3554 ( .IN1(n364), .IN2(\ram[135][6] ), .IN3(n361), .IN4(
        \ram[136][6] ), .Q(n1760) );
  AOI221X1 U3555 ( .IN1(n301), .IN2(\ram[156][6] ), .IN3(n304), .IN4(
        \ram[155][6] ), .IN5(n1761), .QN(n1756) );
  AO22X1 U3556 ( .IN1(n292), .IN2(\ram[159][6] ), .IN3(n289), .IN4(
        \ram[160][6] ), .Q(n1761) );
  AOI221X1 U3557 ( .IN1(n325), .IN2(\ram[148][6] ), .IN3(n328), .IN4(
        \ram[147][6] ), .IN5(n1762), .QN(n1755) );
  AO22X1 U3558 ( .IN1(n316), .IN2(\ram[151][6] ), .IN3(n313), .IN4(
        \ram[152][6] ), .Q(n1762) );
  NAND4X0 U3559 ( .IN1(n1763), .IN2(n1764), .IN3(n1765), .IN4(n1766), .QN(
        n1744) );
  AOI221X1 U3560 ( .IN1(n61), .IN2(\ram[236][6] ), .IN3(n64), .IN4(
        \ram[235][6] ), .IN5(n1767), .QN(n1766) );
  AO22X1 U3561 ( .IN1(n58), .IN2(\ram[237][6] ), .IN3(n55), .IN4(\ram[238][6] ), .Q(n1767) );
  AOI221X1 U3562 ( .IN1(n85), .IN2(\ram[228][6] ), .IN3(n88), .IN4(
        \ram[227][6] ), .IN5(n1768), .QN(n1765) );
  AO22X1 U3563 ( .IN1(n76), .IN2(\ram[231][6] ), .IN3(n73), .IN4(\ram[232][6] ), .Q(n1768) );
  AOI221X1 U3564 ( .IN1(n19), .IN2(\ram[250][6] ), .IN3(n22), .IN4(
        \ram[249][6] ), .IN5(n1769), .QN(n1764) );
  AO22X1 U3565 ( .IN1(n10), .IN2(\ram[253][6] ), .IN3(n7), .IN4(\ram[254][6] ), 
        .Q(n1769) );
  AOI221X1 U3566 ( .IN1(n37), .IN2(\ram[244][6] ), .IN3(n40), .IN4(
        \ram[243][6] ), .IN5(n1770), .QN(n1763) );
  AO22X1 U3567 ( .IN1(n28), .IN2(\ram[247][6] ), .IN3(n25), .IN4(\ram[248][6] ), .Q(n1770) );
  NAND4X0 U3568 ( .IN1(n1771), .IN2(n1772), .IN3(n1773), .IN4(n1774), .QN(
        n1743) );
  AOI221X1 U3569 ( .IN1(n157), .IN2(\ram[204][6] ), .IN3(n160), .IN4(
        \ram[203][6] ), .IN5(n1775), .QN(n1774) );
  AO22X1 U3570 ( .IN1(n148), .IN2(\ram[207][6] ), .IN3(n145), .IN4(
        \ram[208][6] ), .Q(n1775) );
  AOI221X1 U3571 ( .IN1(n181), .IN2(\ram[196][6] ), .IN3(n184), .IN4(
        \ram[195][6] ), .IN5(n1776), .QN(n1773) );
  AO22X1 U3572 ( .IN1(n172), .IN2(\ram[199][6] ), .IN3(n169), .IN4(
        \ram[200][6] ), .Q(n1776) );
  AOI221X1 U3573 ( .IN1(n109), .IN2(\ram[220][6] ), .IN3(n112), .IN4(
        \ram[219][6] ), .IN5(n1777), .QN(n1772) );
  AO22X1 U3574 ( .IN1(n100), .IN2(\ram[223][6] ), .IN3(n97), .IN4(
        \ram[224][6] ), .Q(n1777) );
  AOI221X1 U3575 ( .IN1(n133), .IN2(\ram[212][6] ), .IN3(n136), .IN4(
        \ram[211][6] ), .IN5(n1778), .QN(n1771) );
  AO22X1 U3576 ( .IN1(n124), .IN2(\ram[215][6] ), .IN3(n121), .IN4(
        \ram[216][6] ), .Q(n1778) );
  NAND4X0 U3578 ( .IN1(n1783), .IN2(n1784), .IN3(n1785), .IN4(n1786), .QN(
        n1782) );
  AOI221X1 U3579 ( .IN1(n637), .IN2(\ram[44][6] ), .IN3(n640), .IN4(
        \ram[43][6] ), .IN5(n1787), .QN(n1786) );
  AO22X1 U3580 ( .IN1(n628), .IN2(\ram[47][6] ), .IN3(n625), .IN4(\ram[48][6] ), .Q(n1787) );
  AOI221X1 U3581 ( .IN1(n661), .IN2(\ram[36][6] ), .IN3(n664), .IN4(
        \ram[35][6] ), .IN5(n1788), .QN(n1785) );
  AO22X1 U3582 ( .IN1(n652), .IN2(\ram[39][6] ), .IN3(n649), .IN4(\ram[40][6] ), .Q(n1788) );
  AOI221X1 U3583 ( .IN1(n589), .IN2(\ram[60][6] ), .IN3(n592), .IN4(
        \ram[59][6] ), .IN5(n1789), .QN(n1784) );
  AO22X1 U3584 ( .IN1(n580), .IN2(\ram[63][6] ), .IN3(n577), .IN4(\ram[64][6] ), .Q(n1789) );
  AOI221X1 U3585 ( .IN1(n613), .IN2(\ram[52][6] ), .IN3(n616), .IN4(
        \ram[51][6] ), .IN5(n1790), .QN(n1783) );
  AO22X1 U3586 ( .IN1(n604), .IN2(\ram[55][6] ), .IN3(n601), .IN4(\ram[56][6] ), .Q(n1790) );
  NAND4X0 U3587 ( .IN1(n1791), .IN2(n1792), .IN3(n1793), .IN4(n1794), .QN(
        n1781) );
  AOI221X1 U3588 ( .IN1(n733), .IN2(\ram[12][6] ), .IN3(n736), .IN4(
        \ram[11][6] ), .IN5(n1795), .QN(n1794) );
  AO22X1 U3589 ( .IN1(n724), .IN2(\ram[15][6] ), .IN3(n721), .IN4(\ram[16][6] ), .Q(n1795) );
  AOI221X1 U3590 ( .IN1(n757), .IN2(\ram[4][6] ), .IN3(n760), .IN4(\ram[3][6] ), .IN5(n1796), .QN(n1793) );
  AO22X1 U3591 ( .IN1(n748), .IN2(\ram[7][6] ), .IN3(n745), .IN4(\ram[8][6] ), 
        .Q(n1796) );
  AOI221X1 U3592 ( .IN1(n685), .IN2(\ram[28][6] ), .IN3(n688), .IN4(
        \ram[27][6] ), .IN5(n1797), .QN(n1792) );
  AO22X1 U3593 ( .IN1(n676), .IN2(\ram[31][6] ), .IN3(n673), .IN4(\ram[32][6] ), .Q(n1797) );
  AOI221X1 U3594 ( .IN1(n709), .IN2(\ram[20][6] ), .IN3(n712), .IN4(
        \ram[19][6] ), .IN5(n1798), .QN(n1791) );
  AO22X1 U3595 ( .IN1(n700), .IN2(\ram[23][6] ), .IN3(n697), .IN4(\ram[24][6] ), .Q(n1798) );
  NAND4X0 U3596 ( .IN1(n1799), .IN2(n1800), .IN3(n1801), .IN4(n1802), .QN(
        n1780) );
  AOI221X1 U3597 ( .IN1(n445), .IN2(\ram[108][6] ), .IN3(n448), .IN4(
        \ram[107][6] ), .IN5(n1803), .QN(n1802) );
  AO22X1 U3598 ( .IN1(n436), .IN2(\ram[111][6] ), .IN3(n433), .IN4(
        \ram[112][6] ), .Q(n1803) );
  AOI221X1 U3599 ( .IN1(n469), .IN2(\ram[100][6] ), .IN3(n472), .IN4(
        \ram[99][6] ), .IN5(n1804), .QN(n1801) );
  AO22X1 U3600 ( .IN1(n460), .IN2(\ram[103][6] ), .IN3(n457), .IN4(
        \ram[104][6] ), .Q(n1804) );
  AOI221X1 U3601 ( .IN1(n397), .IN2(\ram[124][6] ), .IN3(n400), .IN4(
        \ram[123][6] ), .IN5(n1805), .QN(n1800) );
  AO22X1 U3602 ( .IN1(n388), .IN2(\ram[127][6] ), .IN3(n385), .IN4(
        \ram[128][6] ), .Q(n1805) );
  AOI221X1 U3603 ( .IN1(n421), .IN2(\ram[116][6] ), .IN3(n424), .IN4(
        \ram[115][6] ), .IN5(n1806), .QN(n1799) );
  AO22X1 U3604 ( .IN1(n412), .IN2(\ram[119][6] ), .IN3(n409), .IN4(
        \ram[120][6] ), .Q(n1806) );
  NAND4X0 U3605 ( .IN1(n1807), .IN2(n1808), .IN3(n1809), .IN4(n1810), .QN(
        n1779) );
  AOI221X1 U3606 ( .IN1(n541), .IN2(\ram[76][6] ), .IN3(n544), .IN4(
        \ram[75][6] ), .IN5(n1811), .QN(n1810) );
  AO22X1 U3607 ( .IN1(n532), .IN2(\ram[79][6] ), .IN3(n529), .IN4(\ram[80][6] ), .Q(n1811) );
  AOI221X1 U3608 ( .IN1(n565), .IN2(\ram[68][6] ), .IN3(n568), .IN4(
        \ram[67][6] ), .IN5(n1812), .QN(n1809) );
  AO22X1 U3609 ( .IN1(n556), .IN2(\ram[71][6] ), .IN3(n553), .IN4(\ram[72][6] ), .Q(n1812) );
  AOI221X1 U3610 ( .IN1(n493), .IN2(\ram[92][6] ), .IN3(n496), .IN4(
        \ram[91][6] ), .IN5(n1813), .QN(n1808) );
  AO22X1 U3611 ( .IN1(n484), .IN2(\ram[95][6] ), .IN3(n481), .IN4(\ram[96][6] ), .Q(n1813) );
  AOI221X1 U3612 ( .IN1(n517), .IN2(\ram[84][6] ), .IN3(n520), .IN4(
        \ram[83][6] ), .IN5(n1814), .QN(n1807) );
  AO22X1 U3613 ( .IN1(n508), .IN2(\ram[87][6] ), .IN3(n505), .IN4(\ram[88][6] ), .Q(n1814) );
  AO22X1 U3614 ( .IN1(n771), .IN2(dataout[7]), .IN3(n4174), .IN4(n1815), .Q(
        n2027) );
  NAND4X0 U3615 ( .IN1(n1816), .IN2(n1817), .IN3(n1818), .IN4(n1819), .QN(
        n1815) );
  NAND4X0 U3617 ( .IN1(n1824), .IN2(n1825), .IN3(n1826), .IN4(n1827), .QN(
        n1823) );
  AOI221X1 U3618 ( .IN1(n259), .IN2(\ram[170][7] ), .IN3(n262), .IN4(
        \ram[169][7] ), .IN5(n1828), .QN(n1827) );
  AO22X1 U3619 ( .IN1(n250), .IN2(\ram[173][7] ), .IN3(n247), .IN4(
        \ram[174][7] ), .Q(n1828) );
  AOI221X1 U3624 ( .IN1(n283), .IN2(\ram[162][7] ), .IN3(n286), .IN4(
        \ram[161][7] ), .IN5(n1834), .QN(n1826) );
  AO22X1 U3625 ( .IN1(n274), .IN2(\ram[165][7] ), .IN3(n271), .IN4(
        \ram[166][7] ), .Q(n1834) );
  AOI221X1 U3630 ( .IN1(n211), .IN2(\ram[186][7] ), .IN3(n214), .IN4(
        \ram[185][7] ), .IN5(n1839), .QN(n1825) );
  AO22X1 U3631 ( .IN1(n196), .IN2(\ram[191][7] ), .IN3(n193), .IN4(
        \ram[192][7] ), .Q(n1839) );
  AOI221X1 U3636 ( .IN1(n235), .IN2(\ram[178][7] ), .IN3(n238), .IN4(
        \ram[177][7] ), .IN5(n1844), .QN(n1824) );
  AO22X1 U3637 ( .IN1(n226), .IN2(\ram[181][7] ), .IN3(n223), .IN4(
        \ram[182][7] ), .Q(n1844) );
  NAND4X0 U3642 ( .IN1(n1845), .IN2(n1846), .IN3(n1847), .IN4(n1848), .QN(
        n1822) );
  AOI221X1 U3643 ( .IN1(n355), .IN2(\ram[138][7] ), .IN3(n358), .IN4(
        \ram[137][7] ), .IN5(n1849), .QN(n1848) );
  AO22X1 U3644 ( .IN1(n346), .IN2(\ram[141][7] ), .IN3(n343), .IN4(
        \ram[142][7] ), .Q(n1849) );
  AOI221X1 U3649 ( .IN1(n379), .IN2(\ram[130][7] ), .IN3(n382), .IN4(
        \ram[129][7] ), .IN5(n1851), .QN(n1847) );
  AO22X1 U3650 ( .IN1(n370), .IN2(\ram[133][7] ), .IN3(n367), .IN4(
        \ram[134][7] ), .Q(n1851) );
  AOI221X1 U3655 ( .IN1(n307), .IN2(\ram[154][7] ), .IN3(n310), .IN4(
        \ram[153][7] ), .IN5(n1852), .QN(n1846) );
  AO22X1 U3656 ( .IN1(n298), .IN2(\ram[157][7] ), .IN3(n295), .IN4(
        \ram[158][7] ), .Q(n1852) );
  AOI221X1 U3661 ( .IN1(n331), .IN2(\ram[146][7] ), .IN3(n334), .IN4(
        \ram[145][7] ), .IN5(n1854), .QN(n1845) );
  AO22X1 U3662 ( .IN1(n322), .IN2(\ram[149][7] ), .IN3(n319), .IN4(
        \ram[150][7] ), .Q(n1854) );
  NAND4X0 U3667 ( .IN1(n1855), .IN2(n1856), .IN3(n1857), .IN4(n1858), .QN(
        n1821) );
  AOI221X1 U3668 ( .IN1(n70), .IN2(\ram[233][7] ), .IN3(n49), .IN4(
        \ram[240][7] ), .IN5(n1859), .QN(n1858) );
  AO22X1 U3669 ( .IN1(n139), .IN2(\ram[210][7] ), .IN3(n52), .IN4(
        \ram[239][7] ), .Q(n1859) );
  AOI221X1 U3674 ( .IN1(n94), .IN2(\ram[225][7] ), .IN3(n79), .IN4(
        \ram[230][7] ), .IN5(n1863), .QN(n1857) );
  AO22X1 U3675 ( .IN1(n67), .IN2(\ram[234][7] ), .IN3(n82), .IN4(\ram[229][7] ), .Q(n1863) );
  AOI221X1 U3680 ( .IN1(n13), .IN2(\ram[252][7] ), .IN3(n16), .IN4(
        \ram[251][7] ), .IN5(n1864), .QN(n1856) );
  AO22X1 U3681 ( .IN1(n91), .IN2(\ram[226][7] ), .IN3(n3), .IN4(\ram[255][7] ), 
        .Q(n1864) );
  AOI221X1 U3686 ( .IN1(n43), .IN2(\ram[242][7] ), .IN3(n46), .IN4(
        \ram[241][7] ), .IN5(n1867), .QN(n1855) );
  AO22X1 U3687 ( .IN1(n34), .IN2(\ram[245][7] ), .IN3(n31), .IN4(\ram[246][7] ), .Q(n1867) );
  NAND4X0 U3692 ( .IN1(n1868), .IN2(n1869), .IN3(n1870), .IN4(n1871), .QN(
        n1820) );
  AOI221X1 U3693 ( .IN1(n166), .IN2(\ram[201][7] ), .IN3(n151), .IN4(
        \ram[206][7] ), .IN5(n1872), .QN(n1871) );
  AO22X1 U3694 ( .IN1(n769), .IN2(\ram[0][7] ), .IN3(n154), .IN4(\ram[205][7] ), .Q(n1872) );
  AOI221X1 U3699 ( .IN1(n190), .IN2(\ram[193][7] ), .IN3(n175), .IN4(
        \ram[198][7] ), .IN5(n1874), .QN(n1870) );
  AO22X1 U3700 ( .IN1(n163), .IN2(\ram[202][7] ), .IN3(n178), .IN4(
        \ram[197][7] ), .Q(n1874) );
  AOI221X1 U3705 ( .IN1(n106), .IN2(\ram[221][7] ), .IN3(n187), .IN4(
        \ram[194][7] ), .IN5(n1875), .QN(n1869) );
  AO22X1 U3706 ( .IN1(n103), .IN2(\ram[222][7] ), .IN3(n118), .IN4(
        \ram[217][7] ), .Q(n1875) );
  AOI221X1 U3711 ( .IN1(n142), .IN2(\ram[209][7] ), .IN3(n127), .IN4(
        \ram[214][7] ), .IN5(n1876), .QN(n1868) );
  AO22X1 U3712 ( .IN1(n115), .IN2(\ram[218][7] ), .IN3(n130), .IN4(
        \ram[213][7] ), .Q(n1876) );
  NAND4X0 U3718 ( .IN1(n1881), .IN2(n1882), .IN3(n1883), .IN4(n1884), .QN(
        n1880) );
  AOI221X1 U3719 ( .IN1(n643), .IN2(\ram[42][7] ), .IN3(n646), .IN4(
        \ram[41][7] ), .IN5(n1885), .QN(n1884) );
  AO22X1 U3720 ( .IN1(n634), .IN2(\ram[45][7] ), .IN3(n631), .IN4(\ram[46][7] ), .Q(n1885) );
  AOI221X1 U3725 ( .IN1(n667), .IN2(\ram[34][7] ), .IN3(n670), .IN4(
        \ram[33][7] ), .IN5(n1887), .QN(n1883) );
  AO22X1 U3726 ( .IN1(n658), .IN2(\ram[37][7] ), .IN3(n655), .IN4(\ram[38][7] ), .Q(n1887) );
  AOI221X1 U3731 ( .IN1(n595), .IN2(\ram[58][7] ), .IN3(n598), .IN4(
        \ram[57][7] ), .IN5(n1888), .QN(n1882) );
  AO22X1 U3732 ( .IN1(n586), .IN2(\ram[61][7] ), .IN3(n583), .IN4(\ram[62][7] ), .Q(n1888) );
  AOI221X1 U3737 ( .IN1(n619), .IN2(\ram[50][7] ), .IN3(n622), .IN4(
        \ram[49][7] ), .IN5(n1890), .QN(n1881) );
  AO22X1 U3738 ( .IN1(n610), .IN2(\ram[53][7] ), .IN3(n607), .IN4(\ram[54][7] ), .Q(n1890) );
  NAND4X0 U3743 ( .IN1(n1891), .IN2(n1892), .IN3(n1893), .IN4(n1894), .QN(
        n1879) );
  AOI221X1 U3744 ( .IN1(n739), .IN2(\ram[10][7] ), .IN3(n742), .IN4(
        \ram[9][7] ), .IN5(n1895), .QN(n1894) );
  AO22X1 U3745 ( .IN1(n730), .IN2(\ram[13][7] ), .IN3(n727), .IN4(\ram[14][7] ), .Q(n1895) );
  AOI221X1 U3750 ( .IN1(n763), .IN2(\ram[2][7] ), .IN3(n766), .IN4(\ram[1][7] ), .IN5(n1896), .QN(n1893) );
  AO22X1 U3751 ( .IN1(n754), .IN2(\ram[5][7] ), .IN3(n751), .IN4(\ram[6][7] ), 
        .Q(n1896) );
  AOI221X1 U3756 ( .IN1(n691), .IN2(\ram[26][7] ), .IN3(n694), .IN4(
        \ram[25][7] ), .IN5(n1897), .QN(n1892) );
  AO22X1 U3757 ( .IN1(n682), .IN2(\ram[29][7] ), .IN3(n679), .IN4(\ram[30][7] ), .Q(n1897) );
  AOI221X1 U3762 ( .IN1(n715), .IN2(\ram[18][7] ), .IN3(n718), .IN4(
        \ram[17][7] ), .IN5(n1899), .QN(n1891) );
  AO22X1 U3763 ( .IN1(n706), .IN2(\ram[21][7] ), .IN3(n703), .IN4(\ram[22][7] ), .Q(n1899) );
  NAND4X0 U3768 ( .IN1(n1900), .IN2(n1901), .IN3(n1902), .IN4(n1903), .QN(
        n1878) );
  AOI221X1 U3769 ( .IN1(n451), .IN2(\ram[106][7] ), .IN3(n454), .IN4(
        \ram[105][7] ), .IN5(n1904), .QN(n1903) );
  AO22X1 U3770 ( .IN1(n442), .IN2(\ram[109][7] ), .IN3(n439), .IN4(
        \ram[110][7] ), .Q(n1904) );
  AOI221X1 U3775 ( .IN1(n475), .IN2(\ram[98][7] ), .IN3(n478), .IN4(
        \ram[97][7] ), .IN5(n1906), .QN(n1902) );
  AO22X1 U3776 ( .IN1(n466), .IN2(\ram[101][7] ), .IN3(n463), .IN4(
        \ram[102][7] ), .Q(n1906) );
  AOI221X1 U3781 ( .IN1(n403), .IN2(\ram[122][7] ), .IN3(n406), .IN4(
        \ram[121][7] ), .IN5(n1907), .QN(n1901) );
  AO22X1 U3782 ( .IN1(n394), .IN2(\ram[125][7] ), .IN3(n391), .IN4(
        \ram[126][7] ), .Q(n1907) );
  AOI221X1 U3787 ( .IN1(n427), .IN2(\ram[114][7] ), .IN3(n430), .IN4(
        \ram[113][7] ), .IN5(n1909), .QN(n1900) );
  AO22X1 U3788 ( .IN1(n418), .IN2(\ram[117][7] ), .IN3(n415), .IN4(
        \ram[118][7] ), .Q(n1909) );
  NAND4X0 U3793 ( .IN1(n1910), .IN2(n1911), .IN3(n1912), .IN4(n1913), .QN(
        n1877) );
  AOI221X1 U3794 ( .IN1(n547), .IN2(\ram[74][7] ), .IN3(n550), .IN4(
        \ram[73][7] ), .IN5(n1914), .QN(n1913) );
  AO22X1 U3795 ( .IN1(n538), .IN2(\ram[77][7] ), .IN3(n535), .IN4(\ram[78][7] ), .Q(n1914) );
  AOI221X1 U3800 ( .IN1(n571), .IN2(\ram[66][7] ), .IN3(n574), .IN4(
        \ram[65][7] ), .IN5(n1916), .QN(n1912) );
  AO22X1 U3801 ( .IN1(n562), .IN2(\ram[69][7] ), .IN3(n559), .IN4(\ram[70][7] ), .Q(n1916) );
  AOI221X1 U3806 ( .IN1(n499), .IN2(\ram[90][7] ), .IN3(n502), .IN4(
        \ram[89][7] ), .IN5(n1917), .QN(n1911) );
  AO22X1 U3807 ( .IN1(n490), .IN2(\ram[93][7] ), .IN3(n487), .IN4(\ram[94][7] ), .Q(n1917) );
  AOI221X1 U3812 ( .IN1(n523), .IN2(\ram[82][7] ), .IN3(n526), .IN4(
        \ram[81][7] ), .IN5(n1919), .QN(n1910) );
  AO22X1 U3813 ( .IN1(n514), .IN2(\ram[85][7] ), .IN3(n511), .IN4(\ram[86][7] ), .Q(n1919) );
  NAND4X0 U3823 ( .IN1(n1930), .IN2(n1931), .IN3(n1932), .IN4(n1933), .QN(
        n1929) );
  AOI221X1 U3824 ( .IN1(n253), .IN2(\ram[172][7] ), .IN3(n256), .IN4(
        \ram[171][7] ), .IN5(n1934), .QN(n1933) );
  AO22X1 U3825 ( .IN1(n244), .IN2(\ram[175][7] ), .IN3(n241), .IN4(
        \ram[176][7] ), .Q(n1934) );
  AOI221X1 U3830 ( .IN1(n277), .IN2(\ram[164][7] ), .IN3(n280), .IN4(
        \ram[163][7] ), .IN5(n1935), .QN(n1932) );
  AO22X1 U3831 ( .IN1(n268), .IN2(\ram[167][7] ), .IN3(n265), .IN4(
        \ram[168][7] ), .Q(n1935) );
  AOI221X1 U3836 ( .IN1(n205), .IN2(\ram[188][7] ), .IN3(n208), .IN4(
        \ram[187][7] ), .IN5(n1940), .QN(n1931) );
  AO22X1 U3837 ( .IN1(n202), .IN2(\ram[189][7] ), .IN3(n199), .IN4(
        \ram[190][7] ), .Q(n1940) );
  AOI221X1 U3842 ( .IN1(n229), .IN2(\ram[180][7] ), .IN3(n232), .IN4(
        \ram[179][7] ), .IN5(n1941), .QN(n1930) );
  AO22X1 U3843 ( .IN1(n220), .IN2(\ram[183][7] ), .IN3(n217), .IN4(
        \ram[184][7] ), .Q(n1941) );
  NAND4X0 U3849 ( .IN1(n1944), .IN2(n1945), .IN3(n1946), .IN4(n1947), .QN(
        n1928) );
  AOI221X1 U3850 ( .IN1(n349), .IN2(\ram[140][7] ), .IN3(n352), .IN4(
        \ram[139][7] ), .IN5(n1948), .QN(n1947) );
  AO22X1 U3851 ( .IN1(n340), .IN2(\ram[143][7] ), .IN3(n337), .IN4(
        \ram[144][7] ), .Q(n1948) );
  AOI221X1 U3856 ( .IN1(n373), .IN2(\ram[132][7] ), .IN3(n376), .IN4(
        \ram[131][7] ), .IN5(n1949), .QN(n1946) );
  AO22X1 U3857 ( .IN1(n364), .IN2(\ram[135][7] ), .IN3(n361), .IN4(
        \ram[136][7] ), .Q(n1949) );
  AOI221X1 U3862 ( .IN1(n301), .IN2(\ram[156][7] ), .IN3(n304), .IN4(
        \ram[155][7] ), .IN5(n1950), .QN(n1945) );
  AO22X1 U3863 ( .IN1(n292), .IN2(\ram[159][7] ), .IN3(n289), .IN4(
        \ram[160][7] ), .Q(n1950) );
  AOI221X1 U3869 ( .IN1(n325), .IN2(\ram[148][7] ), .IN3(n328), .IN4(
        \ram[147][7] ), .IN5(n1952), .QN(n1944) );
  AO22X1 U3870 ( .IN1(n316), .IN2(\ram[151][7] ), .IN3(n313), .IN4(
        \ram[152][7] ), .Q(n1952) );
  NAND4X0 U3876 ( .IN1(n1954), .IN2(n1955), .IN3(n1956), .IN4(n1957), .QN(
        n1927) );
  AOI221X1 U3877 ( .IN1(n61), .IN2(\ram[236][7] ), .IN3(n64), .IN4(
        \ram[235][7] ), .IN5(n1958), .QN(n1957) );
  AO22X1 U3878 ( .IN1(n58), .IN2(\ram[237][7] ), .IN3(n55), .IN4(\ram[238][7] ), .Q(n1958) );
  AOI221X1 U3883 ( .IN1(n85), .IN2(\ram[228][7] ), .IN3(n88), .IN4(
        \ram[227][7] ), .IN5(n1959), .QN(n1956) );
  AO22X1 U3884 ( .IN1(n76), .IN2(\ram[231][7] ), .IN3(n73), .IN4(\ram[232][7] ), .Q(n1959) );
  AOI221X1 U3889 ( .IN1(n19), .IN2(\ram[250][7] ), .IN3(n22), .IN4(
        \ram[249][7] ), .IN5(n1960), .QN(n1955) );
  AO22X1 U3890 ( .IN1(n10), .IN2(\ram[253][7] ), .IN3(n7), .IN4(\ram[254][7] ), 
        .Q(n1960) );
  AOI221X1 U3899 ( .IN1(n37), .IN2(\ram[244][7] ), .IN3(n40), .IN4(
        \ram[243][7] ), .IN5(n1963), .QN(n1954) );
  AO22X1 U3900 ( .IN1(n28), .IN2(\ram[247][7] ), .IN3(n25), .IN4(\ram[248][7] ), .Q(n1963) );
  NAND4X0 U3906 ( .IN1(n1965), .IN2(n1966), .IN3(n1967), .IN4(n1968), .QN(
        n1926) );
  AOI221X1 U3907 ( .IN1(n157), .IN2(\ram[204][7] ), .IN3(n160), .IN4(
        \ram[203][7] ), .IN5(n1969), .QN(n1968) );
  AO22X1 U3908 ( .IN1(n148), .IN2(\ram[207][7] ), .IN3(n145), .IN4(
        \ram[208][7] ), .Q(n1969) );
  AOI221X1 U3913 ( .IN1(n181), .IN2(\ram[196][7] ), .IN3(n184), .IN4(
        \ram[195][7] ), .IN5(n1970), .QN(n1967) );
  AO22X1 U3914 ( .IN1(n172), .IN2(\ram[199][7] ), .IN3(n169), .IN4(
        \ram[200][7] ), .Q(n1970) );
  AOI221X1 U3920 ( .IN1(n109), .IN2(\ram[220][7] ), .IN3(n112), .IN4(
        \ram[219][7] ), .IN5(n1972), .QN(n1966) );
  AO22X1 U3921 ( .IN1(n100), .IN2(\ram[223][7] ), .IN3(n97), .IN4(
        \ram[224][7] ), .Q(n1972) );
  AOI221X1 U3927 ( .IN1(n133), .IN2(\ram[212][7] ), .IN3(n136), .IN4(
        \ram[211][7] ), .IN5(n1973), .QN(n1965) );
  AO22X1 U3928 ( .IN1(n124), .IN2(\ram[215][7] ), .IN3(n121), .IN4(
        \ram[216][7] ), .Q(n1973) );
  NAND4X0 U3936 ( .IN1(n1980), .IN2(n1981), .IN3(n1982), .IN4(n1983), .QN(
        n1979) );
  AOI221X1 U3937 ( .IN1(n637), .IN2(\ram[44][7] ), .IN3(n640), .IN4(
        \ram[43][7] ), .IN5(n1984), .QN(n1983) );
  AO22X1 U3938 ( .IN1(n628), .IN2(\ram[47][7] ), .IN3(n625), .IN4(\ram[48][7] ), .Q(n1984) );
  AOI221X1 U3943 ( .IN1(n661), .IN2(\ram[36][7] ), .IN3(n664), .IN4(
        \ram[35][7] ), .IN5(n1985), .QN(n1982) );
  AO22X1 U3944 ( .IN1(n652), .IN2(\ram[39][7] ), .IN3(n649), .IN4(\ram[40][7] ), .Q(n1985) );
  AOI221X1 U3949 ( .IN1(n589), .IN2(\ram[60][7] ), .IN3(n592), .IN4(
        \ram[59][7] ), .IN5(n1986), .QN(n1981) );
  AO22X1 U3950 ( .IN1(n580), .IN2(\ram[63][7] ), .IN3(n577), .IN4(\ram[64][7] ), .Q(n1986) );
  AOI221X1 U3955 ( .IN1(n613), .IN2(\ram[52][7] ), .IN3(n616), .IN4(
        \ram[51][7] ), .IN5(n1987), .QN(n1980) );
  AO22X1 U3956 ( .IN1(n604), .IN2(\ram[55][7] ), .IN3(n601), .IN4(\ram[56][7] ), .Q(n1987) );
  NAND4X0 U3962 ( .IN1(n1989), .IN2(n1990), .IN3(n1991), .IN4(n1992), .QN(
        n1978) );
  AOI221X1 U3963 ( .IN1(n733), .IN2(\ram[12][7] ), .IN3(n736), .IN4(
        \ram[11][7] ), .IN5(n1993), .QN(n1992) );
  AO22X1 U3964 ( .IN1(n724), .IN2(\ram[15][7] ), .IN3(n721), .IN4(\ram[16][7] ), .Q(n1993) );
  AOI221X1 U3969 ( .IN1(n757), .IN2(\ram[4][7] ), .IN3(n760), .IN4(\ram[3][7] ), .IN5(n1994), .QN(n1991) );
  AO22X1 U3970 ( .IN1(n748), .IN2(\ram[7][7] ), .IN3(n745), .IN4(\ram[8][7] ), 
        .Q(n1994) );
  AOI221X1 U3976 ( .IN1(n685), .IN2(\ram[28][7] ), .IN3(n688), .IN4(
        \ram[27][7] ), .IN5(n1995), .QN(n1990) );
  AO22X1 U3977 ( .IN1(n676), .IN2(\ram[31][7] ), .IN3(n673), .IN4(\ram[32][7] ), .Q(n1995) );
  AOI221X1 U3983 ( .IN1(n709), .IN2(\ram[20][7] ), .IN3(n712), .IN4(
        \ram[19][7] ), .IN5(n1996), .QN(n1989) );
  AO22X1 U3984 ( .IN1(n700), .IN2(\ram[23][7] ), .IN3(n697), .IN4(\ram[24][7] ), .Q(n1996) );
  NAND4X0 U3991 ( .IN1(n1997), .IN2(n1998), .IN3(n1999), .IN4(n2000), .QN(
        n1977) );
  AOI221X1 U3992 ( .IN1(n445), .IN2(\ram[108][7] ), .IN3(n448), .IN4(
        \ram[107][7] ), .IN5(n2001), .QN(n2000) );
  AO22X1 U3993 ( .IN1(n436), .IN2(\ram[111][7] ), .IN3(n433), .IN4(
        \ram[112][7] ), .Q(n2001) );
  AOI221X1 U3998 ( .IN1(n469), .IN2(\ram[100][7] ), .IN3(n472), .IN4(
        \ram[99][7] ), .IN5(n2002), .QN(n1999) );
  AO22X1 U3999 ( .IN1(n460), .IN2(\ram[103][7] ), .IN3(n457), .IN4(
        \ram[104][7] ), .Q(n2002) );
  AOI221X1 U4004 ( .IN1(n397), .IN2(\ram[124][7] ), .IN3(n400), .IN4(
        \ram[123][7] ), .IN5(n2003), .QN(n1998) );
  AO22X1 U4005 ( .IN1(n388), .IN2(\ram[127][7] ), .IN3(n385), .IN4(
        \ram[128][7] ), .Q(n2003) );
  AOI221X1 U4013 ( .IN1(n421), .IN2(\ram[116][7] ), .IN3(n424), .IN4(
        \ram[115][7] ), .IN5(n2004), .QN(n1997) );
  AO22X1 U4014 ( .IN1(n412), .IN2(\ram[119][7] ), .IN3(n409), .IN4(
        \ram[120][7] ), .Q(n2004) );
  NAND4X0 U4021 ( .IN1(n2008), .IN2(n2009), .IN3(n2010), .IN4(n2011), .QN(
        n1976) );
  AOI221X1 U4022 ( .IN1(n541), .IN2(\ram[76][7] ), .IN3(n544), .IN4(
        \ram[75][7] ), .IN5(n2012), .QN(n2011) );
  AO22X1 U4023 ( .IN1(n532), .IN2(\ram[79][7] ), .IN3(n529), .IN4(\ram[80][7] ), .Q(n2012) );
  AOI221X1 U4028 ( .IN1(n565), .IN2(\ram[68][7] ), .IN3(n568), .IN4(
        \ram[67][7] ), .IN5(n2013), .QN(n2010) );
  AO22X1 U4029 ( .IN1(n556), .IN2(\ram[71][7] ), .IN3(n553), .IN4(\ram[72][7] ), .Q(n2013) );
  AOI221X1 U4036 ( .IN1(n493), .IN2(\ram[92][7] ), .IN3(n496), .IN4(
        \ram[91][7] ), .IN5(n2014), .QN(n2009) );
  AO22X1 U4037 ( .IN1(n484), .IN2(\ram[95][7] ), .IN3(n481), .IN4(\ram[96][7] ), .Q(n2014) );
  AOI221X1 U4050 ( .IN1(n517), .IN2(\ram[84][7] ), .IN3(n520), .IN4(
        \ram[83][7] ), .IN5(n2017), .QN(n2008) );
  AO22X1 U4051 ( .IN1(n508), .IN2(\ram[87][7] ), .IN3(n505), .IN4(\ram[88][7] ), .Q(n2017) );
  INVX0 U11 ( .IN(W), .QN(n4175) );
  INVX0 U12 ( .IN(n1), .QN(n387) );
  NAND2X0 U21 ( .IN1(n3), .IN2(n4), .QN(n1) );
  INVX0 U22 ( .IN(n11), .QN(n2006) );
  INVX0 U31 ( .IN(n17), .QN(n2007) );
  INVX0 U32 ( .IN(n35), .QN(n4113) );
  INVX0 U41 ( .IN(n41), .QN(n4144) );
  INVX0 U42 ( .IN(n59), .QN(n765) );
  INVX0 U51 ( .IN(n68), .QN(n429) );
  INVX0 U52 ( .IN(n83), .QN(n4114) );
  INVX0 U61 ( .IN(n92), .QN(n621) );
  INVX0 U62 ( .IN(n104), .QN(n477) );
  INVX0 U71 ( .IN(n107), .QN(n759) );
  INVX0 U72 ( .IN(n131), .QN(n4111) );
  INVX0 U81 ( .IN(n140), .QN(n612) );
  INVX0 U82 ( .IN(n155), .QN(n762) );
  INVX0 U91 ( .IN(n164), .QN(n426) );
  INVX0 U92 ( .IN(n179), .QN(n4112) );
  INVX0 U101 ( .IN(n188), .QN(n615) );
  INVX0 U102 ( .IN(n203), .QN(n1974) );
  INVX0 U111 ( .IN(n209), .QN(n4085) );
  INVX0 U112 ( .IN(n227), .QN(n4117) );
  INVX0 U121 ( .IN(n233), .QN(n4149) );
  INVX0 U122 ( .IN(n251), .QN(n1975) );
  INVX0 U131 ( .IN(n257), .QN(n4086) );
  INVX0 U132 ( .IN(n275), .QN(n4118) );
  INVX0 U141 ( .IN(n281), .QN(n4150) );
  INVX0 U142 ( .IN(n299), .QN(n768) );
  INVX0 U151 ( .IN(n305), .QN(n4083) );
  INVX0 U152 ( .IN(n323), .QN(n4115) );
  INVX0 U161 ( .IN(n329), .QN(n4147) );
  INVX0 U162 ( .IN(n347), .QN(n770) );
  INVX0 U171 ( .IN(n353), .QN(n4084) );
  INVX0 U172 ( .IN(n371), .QN(n4116) );
  INVX0 U181 ( .IN(n377), .QN(n4148) );
  INVX0 U182 ( .IN(n395), .QN(n741) );
  INVX0 U191 ( .IN(n401), .QN(n2018) );
  INVX0 U192 ( .IN(n419), .QN(n4105) );
  INVX0 U201 ( .IN(n425), .QN(n4137) );
  INVX0 U202 ( .IN(n443), .QN(n744) );
  INVX0 U211 ( .IN(n449), .QN(n2019) );
  INVX0 U212 ( .IN(n467), .QN(n4106) );
  INVX0 U221 ( .IN(n473), .QN(n4138) );
  INVX0 U222 ( .IN(n491), .QN(n735) );
  INVX0 U231 ( .IN(n497), .QN(n2015) );
  INVX0 U232 ( .IN(n515), .QN(n4103) );
  INVX0 U241 ( .IN(n521), .QN(n4135) );
  INVX0 U242 ( .IN(n539), .QN(n738) );
  INVX0 U251 ( .IN(n545), .QN(n2016) );
  INVX0 U252 ( .IN(n563), .QN(n4104) );
  INVX0 U261 ( .IN(n569), .QN(n4136) );
  INVX0 U262 ( .IN(n587), .QN(n753) );
  INVX0 U271 ( .IN(n593), .QN(n4078) );
  INVX0 U272 ( .IN(n611), .QN(n4109) );
  INVX0 U281 ( .IN(n617), .QN(n4141) );
  INVX0 U282 ( .IN(n635), .QN(n756) );
  INVX0 U291 ( .IN(n641), .QN(n4079) );
  INVX0 U292 ( .IN(n659), .QN(n4110) );
  INVX0 U301 ( .IN(n665), .QN(n4142) );
  INVX0 U302 ( .IN(n683), .QN(n747) );
  INVX0 U311 ( .IN(n689), .QN(n4076) );
  INVX0 U312 ( .IN(n707), .QN(n4107) );
  INVX0 U321 ( .IN(n713), .QN(n4139) );
  INVX0 U322 ( .IN(n731), .QN(n750) );
  INVX0 U331 ( .IN(n737), .QN(n4077) );
  INVX0 U332 ( .IN(n755), .QN(n4108) );
  INVX0 U341 ( .IN(n761), .QN(n4140) );
  INVX0 U342 ( .IN(n8), .QN(n444) );
  INVX0 U351 ( .IN(n26), .QN(n570) );
  INVX0 U352 ( .IN(n32), .QN(n666) );
  INVX0 U361 ( .IN(n56), .QN(n447) );
  INVX0 U362 ( .IN(n65), .QN(n4082) );
  INVX0 U371 ( .IN(n74), .QN(n573) );
  INVX0 U372 ( .IN(n89), .QN(n4145) );
  INVX0 U381 ( .IN(n98), .QN(n372) );
  INVX0 U382 ( .IN(n101), .QN(n4098) );
  INVX0 U391 ( .IN(n113), .QN(n4080) );
  INVX0 U392 ( .IN(n122), .QN(n564) );
  INVX0 U401 ( .IN(n137), .QN(n4146) );
  INVX0 U402 ( .IN(n146), .QN(n375) );
  INVX0 U411 ( .IN(n161), .QN(n4081) );
  INVX0 U412 ( .IN(n170), .QN(n567) );
  INVX0 U421 ( .IN(n194), .QN(n393) );
  INVX0 U422 ( .IN(n200), .QN(n450) );
  INVX0 U431 ( .IN(n218), .QN(n582) );
  INVX0 U432 ( .IN(n224), .QN(n678) );
  INVX0 U441 ( .IN(n242), .QN(n384) );
  INVX0 U442 ( .IN(n248), .QN(n489) );
  INVX0 U451 ( .IN(n266), .QN(n585) );
  INVX0 U452 ( .IN(n272), .QN(n681) );
  INVX0 U461 ( .IN(n290), .QN(n378) );
  INVX0 U462 ( .IN(n296), .QN(n483) );
  INVX0 U471 ( .IN(n314), .QN(n576) );
  INVX0 U472 ( .IN(n320), .QN(n672) );
  INVX0 U481 ( .IN(n338), .QN(n381) );
  INVX0 U482 ( .IN(n344), .QN(n486) );
  INVX0 U491 ( .IN(n362), .QN(n579) );
  INVX0 U492 ( .IN(n368), .QN(n675) );
  INVX0 U501 ( .IN(n386), .QN(n354) );
  INVX0 U502 ( .IN(n392), .QN(n459) );
  INVX0 U511 ( .IN(n410), .QN(n546) );
  INVX0 U512 ( .IN(n416), .QN(n642) );
  INVX0 U521 ( .IN(n434), .QN(n357) );
  INVX0 U522 ( .IN(n440), .QN(n462) );
  INVX0 U531 ( .IN(n458), .QN(n549) );
  INVX0 U532 ( .IN(n464), .QN(n645) );
  INVX0 U541 ( .IN(n482), .QN(n348) );
  INVX0 U542 ( .IN(n488), .QN(n453) );
  INVX0 U551 ( .IN(n506), .QN(n540) );
  INVX0 U552 ( .IN(n512), .QN(n636) );
  INVX0 U561 ( .IN(n530), .QN(n351) );
  INVX0 U562 ( .IN(n536), .QN(n456) );
  INVX0 U571 ( .IN(n554), .QN(n543) );
  INVX0 U572 ( .IN(n560), .QN(n639) );
  INVX0 U581 ( .IN(n578), .QN(n366) );
  INVX0 U582 ( .IN(n584), .QN(n471) );
  INVX0 U591 ( .IN(n602), .QN(n558) );
  INVX0 U592 ( .IN(n608), .QN(n654) );
  INVX0 U601 ( .IN(n626), .QN(n369) );
  INVX0 U602 ( .IN(n632), .QN(n474) );
  INVX0 U611 ( .IN(n650), .QN(n561) );
  INVX0 U612 ( .IN(n656), .QN(n657) );
  INVX0 U621 ( .IN(n674), .QN(n360) );
  INVX0 U622 ( .IN(n680), .QN(n465) );
  INVX0 U631 ( .IN(n698), .QN(n552) );
  INVX0 U632 ( .IN(n704), .QN(n648) );
  INVX0 U641 ( .IN(n722), .QN(n363) );
  INVX0 U642 ( .IN(n728), .QN(n468) );
  INVX0 U651 ( .IN(n746), .QN(n555) );
  INVX0 U652 ( .IN(n752), .QN(n651) );
  INVX0 U661 ( .IN(n767), .QN(n4132) );
  INVX0 U662 ( .IN(n5), .QN(n4087) );
  INVX0 U671 ( .IN(n23), .QN(n717) );
  INVX0 U672 ( .IN(n29), .QN(n4161) );
  INVX0 U681 ( .IN(n50), .QN(n390) );
  INVX0 U682 ( .IN(n53), .QN(n4088) );
  INVX0 U691 ( .IN(n71), .QN(n720) );
  INVX0 U692 ( .IN(n80), .QN(n669) );
  INVX0 U701 ( .IN(n95), .QN(n4127) );
  INVX0 U702 ( .IN(n116), .QN(n423) );
  INVX0 U711 ( .IN(n119), .QN(n711) );
  INVX0 U712 ( .IN(n128), .QN(n660) );
  INVX0 U721 ( .IN(n143), .QN(n4128) );
  INVX0 U722 ( .IN(n152), .QN(n480) );
  INVX0 U731 ( .IN(n167), .QN(n714) );
  INVX0 U732 ( .IN(n176), .QN(n663) );
  INVX0 U741 ( .IN(n191), .QN(n4134) );
  INVX0 U742 ( .IN(n197), .QN(n4089) );
  INVX0 U751 ( .IN(n215), .QN(n729) );
  INVX0 U752 ( .IN(n221), .QN(n4165) );
  INVX0 U761 ( .IN(n239), .QN(n4131) );
  INVX0 U762 ( .IN(n245), .QN(n4102) );
  INVX0 U771 ( .IN(n263), .QN(n732) );
  INVX0 U772 ( .IN(n269), .QN(n4166) );
  INVX0 U781 ( .IN(n287), .QN(n4129) );
  INVX0 U782 ( .IN(n293), .QN(n4100) );
  INVX0 U791 ( .IN(n311), .QN(n723) );
  INVX0 U792 ( .IN(n317), .QN(n4163) );
  INVX0 U801 ( .IN(n335), .QN(n4130) );
  INVX0 U802 ( .IN(n341), .QN(n4101) );
  INVX0 U811 ( .IN(n359), .QN(n726) );
  INVX0 U812 ( .IN(n365), .QN(n4164) );
  INVX0 U821 ( .IN(n383), .QN(n4121) );
  INVX0 U822 ( .IN(n389), .QN(n4092) );
  INVX0 U831 ( .IN(n407), .QN(n693) );
  INVX0 U832 ( .IN(n413), .QN(n4153) );
  INVX0 U841 ( .IN(n431), .QN(n4122) );
  INVX0 U842 ( .IN(n437), .QN(n4093) );
  INVX0 U851 ( .IN(n455), .QN(n696) );
  INVX0 U852 ( .IN(n461), .QN(n4154) );
  INVX0 U861 ( .IN(n479), .QN(n4119) );
  INVX0 U862 ( .IN(n485), .QN(n4090) );
  INVX0 U871 ( .IN(n503), .QN(n687) );
  INVX0 U872 ( .IN(n509), .QN(n4151) );
  INVX0 U881 ( .IN(n527), .QN(n4120) );
  INVX0 U882 ( .IN(n533), .QN(n4091) );
  INVX0 U891 ( .IN(n551), .QN(n690) );
  INVX0 U892 ( .IN(n557), .QN(n4152) );
  INVX0 U901 ( .IN(n575), .QN(n4125) );
  INVX0 U902 ( .IN(n581), .QN(n4096) );
  INVX0 U911 ( .IN(n599), .QN(n705) );
  INVX0 U912 ( .IN(n605), .QN(n4157) );
  INVX0 U921 ( .IN(n623), .QN(n4126) );
  INVX0 U922 ( .IN(n629), .QN(n4097) );
  INVX0 U931 ( .IN(n647), .QN(n708) );
  INVX0 U932 ( .IN(n653), .QN(n4158) );
  INVX0 U941 ( .IN(n671), .QN(n4123) );
  INVX0 U942 ( .IN(n677), .QN(n4094) );
  INVX0 U951 ( .IN(n695), .QN(n699) );
  INVX0 U952 ( .IN(n701), .QN(n4155) );
  INVX0 U961 ( .IN(n719), .QN(n4124) );
  INVX0 U962 ( .IN(n725), .QN(n4095) );
  INVX0 U971 ( .IN(n743), .QN(n702) );
  INVX0 U972 ( .IN(n749), .QN(n4156) );
  INVX0 U981 ( .IN(n14), .QN(n345) );
  INVX0 U982 ( .IN(n20), .QN(n396) );
  INVX0 U991 ( .IN(n38), .QN(n522) );
  INVX0 U992 ( .IN(n44), .QN(n618) );
  INVX0 U1001 ( .IN(n47), .QN(n4133) );
  INVX0 U1002 ( .IN(n62), .QN(n330) );
  INVX0 U1011 ( .IN(n77), .QN(n4162) );
  INVX0 U1012 ( .IN(n86), .QN(n525) );
  INVX0 U1021 ( .IN(n110), .QN(n324) );
  INVX0 U1022 ( .IN(n125), .QN(n4159) );
  INVX0 U1031 ( .IN(n134), .QN(n516) );
  INVX0 U1032 ( .IN(n149), .QN(n4099) );
  INVX0 U1041 ( .IN(n158), .QN(n327) );
  INVX0 U1042 ( .IN(n173), .QN(n4160) );
  INVX0 U1051 ( .IN(n182), .QN(n519) );
  INVX0 U1052 ( .IN(n185), .QN(n4143) );
  INVX0 U1061 ( .IN(n206), .QN(n339) );
  INVX0 U1062 ( .IN(n212), .QN(n438) );
  INVX0 U1071 ( .IN(n230), .QN(n534) );
  INVX0 U1072 ( .IN(n236), .QN(n630) );
  INVX0 U1081 ( .IN(n254), .QN(n342) );
  INVX0 U1082 ( .IN(n260), .QN(n441) );
  INVX0 U1091 ( .IN(n278), .QN(n537) );
  INVX0 U1092 ( .IN(n284), .QN(n633) );
  INVX0 U1101 ( .IN(n302), .QN(n333) );
  INVX0 U1102 ( .IN(n308), .QN(n432) );
  INVX0 U1111 ( .IN(n326), .QN(n528) );
  INVX0 U1112 ( .IN(n332), .QN(n624) );
  INVX0 U1121 ( .IN(n350), .QN(n336) );
  INVX0 U1122 ( .IN(n356), .QN(n435) );
  INVX0 U1131 ( .IN(n374), .QN(n531) );
  INVX0 U1132 ( .IN(n380), .QN(n627) );
  INVX0 U1141 ( .IN(n398), .QN(n306) );
  INVX0 U1142 ( .IN(n404), .QN(n405) );
  INVX0 U1151 ( .IN(n422), .QN(n498) );
  INVX0 U1152 ( .IN(n428), .QN(n594) );
  INVX0 U1161 ( .IN(n446), .QN(n309) );
  INVX0 U1162 ( .IN(n452), .QN(n408) );
  INVX0 U1171 ( .IN(n470), .QN(n501) );
  INVX0 U1172 ( .IN(n476), .QN(n597) );
  INVX0 U1181 ( .IN(n494), .QN(n300) );
  INVX0 U1182 ( .IN(n500), .QN(n399) );
  INVX0 U1191 ( .IN(n518), .QN(n492) );
  INVX0 U1192 ( .IN(n524), .QN(n588) );
  INVX0 U1201 ( .IN(n542), .QN(n303) );
  INVX0 U1202 ( .IN(n548), .QN(n402) );
  INVX0 U1211 ( .IN(n566), .QN(n495) );
  INVX0 U1212 ( .IN(n572), .QN(n591) );
  INVX0 U1221 ( .IN(n590), .QN(n318) );
  INVX0 U1222 ( .IN(n596), .QN(n417) );
  INVX0 U1231 ( .IN(n614), .QN(n510) );
  INVX0 U1232 ( .IN(n620), .QN(n606) );
  INVX0 U1241 ( .IN(n638), .QN(n321) );
  INVX0 U1242 ( .IN(n644), .QN(n420) );
  INVX0 U1251 ( .IN(n662), .QN(n513) );
  INVX0 U1252 ( .IN(n668), .QN(n609) );
  INVX0 U1261 ( .IN(n686), .QN(n312) );
  INVX0 U1262 ( .IN(n692), .QN(n411) );
  INVX0 U1271 ( .IN(n710), .QN(n504) );
  INVX0 U1272 ( .IN(n716), .QN(n600) );
  INVX0 U1281 ( .IN(n734), .QN(n315) );
  INVX0 U1282 ( .IN(n740), .QN(n414) );
  INVX0 U1291 ( .IN(n758), .QN(n507) );
  INVX0 U1292 ( .IN(n764), .QN(n603) );
  INVX0 U1301 ( .IN(n33), .QN(n30) );
  INVX0 U1302 ( .IN(n33), .QN(n27) );
  INVX0 U1311 ( .IN(n33), .QN(n24) );
  INVX0 U1312 ( .IN(n33), .QN(n21) );
  INVX0 U1321 ( .IN(n33), .QN(n18) );
  INVX0 U1322 ( .IN(n33), .QN(n15) );
  INVX0 U1331 ( .IN(n33), .QN(n12) );
  INVX0 U1332 ( .IN(n33), .QN(n9) );
  INVX0 U1341 ( .IN(n33), .QN(n6) );
  INVX0 U1342 ( .IN(n33), .QN(n2) );
  NAND2X0 U1351 ( .IN1(n16), .IN2(n30), .QN(n14) );
  NAND2X0 U1352 ( .IN1(n19), .IN2(n30), .QN(n17) );
  NAND2X0 U1361 ( .IN1(n22), .IN2(n30), .QN(n20) );
  NAND2X0 U1362 ( .IN1(n25), .IN2(n30), .QN(n23) );
  NAND2X0 U1371 ( .IN1(n28), .IN2(n30), .QN(n26) );
  NAND2X0 U1372 ( .IN1(n31), .IN2(n30), .QN(n29) );
  NAND2X0 U1381 ( .IN1(n34), .IN2(n30), .QN(n32) );
  NAND2X0 U1382 ( .IN1(n37), .IN2(n30), .QN(n35) );
  NAND2X0 U1391 ( .IN1(n40), .IN2(n30), .QN(n38) );
  NAND2X0 U1392 ( .IN1(n43), .IN2(n30), .QN(n41) );
  NAND2X0 U1401 ( .IN1(n46), .IN2(n30), .QN(n44) );
  NAND2X0 U1402 ( .IN1(n49), .IN2(n30), .QN(n47) );
  NAND2X0 U1411 ( .IN1(n52), .IN2(n27), .QN(n50) );
  NAND2X0 U1412 ( .IN1(n55), .IN2(n27), .QN(n53) );
  NAND2X0 U1421 ( .IN1(n58), .IN2(n27), .QN(n56) );
  NAND2X0 U1422 ( .IN1(n61), .IN2(n27), .QN(n59) );
  NAND2X0 U1431 ( .IN1(n64), .IN2(n27), .QN(n62) );
  NAND2X0 U1432 ( .IN1(n67), .IN2(n27), .QN(n65) );
  NAND2X0 U1441 ( .IN1(n70), .IN2(n27), .QN(n68) );
  NAND2X0 U1442 ( .IN1(n73), .IN2(n27), .QN(n71) );
  NAND2X0 U1451 ( .IN1(n76), .IN2(n27), .QN(n74) );
  NAND2X0 U1452 ( .IN1(n79), .IN2(n27), .QN(n77) );
  NAND2X0 U1461 ( .IN1(n82), .IN2(n27), .QN(n80) );
  NAND2X0 U1462 ( .IN1(n85), .IN2(n27), .QN(n83) );
  NAND2X0 U1471 ( .IN1(n88), .IN2(n24), .QN(n86) );
  NAND2X0 U1472 ( .IN1(n91), .IN2(n24), .QN(n89) );
  NAND2X0 U1481 ( .IN1(n94), .IN2(n24), .QN(n92) );
  NAND2X0 U1482 ( .IN1(n97), .IN2(n24), .QN(n95) );
  NAND2X0 U1491 ( .IN1(n100), .IN2(n24), .QN(n98) );
  NAND2X0 U1492 ( .IN1(n103), .IN2(n24), .QN(n101) );
  NAND2X0 U1501 ( .IN1(n106), .IN2(n24), .QN(n104) );
  NAND2X0 U1502 ( .IN1(n109), .IN2(n24), .QN(n107) );
  NAND2X0 U1511 ( .IN1(n112), .IN2(n24), .QN(n110) );
  NAND2X0 U1512 ( .IN1(n115), .IN2(n24), .QN(n113) );
  NAND2X0 U1521 ( .IN1(n118), .IN2(n24), .QN(n116) );
  NAND2X0 U1522 ( .IN1(n121), .IN2(n24), .QN(n119) );
  NAND2X0 U1531 ( .IN1(n124), .IN2(n21), .QN(n122) );
  NAND2X0 U1532 ( .IN1(n127), .IN2(n21), .QN(n125) );
  NAND2X0 U1541 ( .IN1(n130), .IN2(n21), .QN(n128) );
  NAND2X0 U1542 ( .IN1(n133), .IN2(n21), .QN(n131) );
  NAND2X0 U1551 ( .IN1(n136), .IN2(n21), .QN(n134) );
  NAND2X0 U1552 ( .IN1(n139), .IN2(n21), .QN(n137) );
  NAND2X0 U1561 ( .IN1(n142), .IN2(n21), .QN(n140) );
  NAND2X0 U1562 ( .IN1(n145), .IN2(n21), .QN(n143) );
  NAND2X0 U1571 ( .IN1(n148), .IN2(n21), .QN(n146) );
  NAND2X0 U1572 ( .IN1(n151), .IN2(n21), .QN(n149) );
  NAND2X0 U1581 ( .IN1(n154), .IN2(n21), .QN(n152) );
  NAND2X0 U1582 ( .IN1(n157), .IN2(n21), .QN(n155) );
  NAND2X0 U1591 ( .IN1(n160), .IN2(n18), .QN(n158) );
  NAND2X0 U1592 ( .IN1(n163), .IN2(n18), .QN(n161) );
  NAND2X0 U1601 ( .IN1(n166), .IN2(n18), .QN(n164) );
  NAND2X0 U1602 ( .IN1(n169), .IN2(n18), .QN(n167) );
  NAND2X0 U1611 ( .IN1(n172), .IN2(n18), .QN(n170) );
  NAND2X0 U1612 ( .IN1(n175), .IN2(n18), .QN(n173) );
  NAND2X0 U1621 ( .IN1(n178), .IN2(n18), .QN(n176) );
  NAND2X0 U1622 ( .IN1(n181), .IN2(n18), .QN(n179) );
  NAND2X0 U1631 ( .IN1(n184), .IN2(n18), .QN(n182) );
  NAND2X0 U1632 ( .IN1(n187), .IN2(n18), .QN(n185) );
  NAND2X0 U1641 ( .IN1(n190), .IN2(n18), .QN(n188) );
  NAND2X0 U1642 ( .IN1(n193), .IN2(n18), .QN(n191) );
  NAND2X0 U1651 ( .IN1(n196), .IN2(n15), .QN(n194) );
  NAND2X0 U1652 ( .IN1(n199), .IN2(n15), .QN(n197) );
  NAND2X0 U1661 ( .IN1(n202), .IN2(n15), .QN(n200) );
  NAND2X0 U1662 ( .IN1(n205), .IN2(n15), .QN(n203) );
  NAND2X0 U1671 ( .IN1(n208), .IN2(n15), .QN(n206) );
  NAND2X0 U1672 ( .IN1(n211), .IN2(n15), .QN(n209) );
  NAND2X0 U1681 ( .IN1(n214), .IN2(n15), .QN(n212) );
  NAND2X0 U1682 ( .IN1(n217), .IN2(n15), .QN(n215) );
  NAND2X0 U1691 ( .IN1(n220), .IN2(n15), .QN(n218) );
  NAND2X0 U1692 ( .IN1(n223), .IN2(n15), .QN(n221) );
  NAND2X0 U1701 ( .IN1(n226), .IN2(n15), .QN(n224) );
  NAND2X0 U1702 ( .IN1(n229), .IN2(n15), .QN(n227) );
  NAND2X0 U1711 ( .IN1(n232), .IN2(n12), .QN(n230) );
  NAND2X0 U1712 ( .IN1(n235), .IN2(n12), .QN(n233) );
  NAND2X0 U1721 ( .IN1(n238), .IN2(n12), .QN(n236) );
  NAND2X0 U1722 ( .IN1(n241), .IN2(n12), .QN(n239) );
  NAND2X0 U1731 ( .IN1(n244), .IN2(n12), .QN(n242) );
  NAND2X0 U1732 ( .IN1(n247), .IN2(n12), .QN(n245) );
  NAND2X0 U1741 ( .IN1(n250), .IN2(n12), .QN(n248) );
  NAND2X0 U1742 ( .IN1(n253), .IN2(n12), .QN(n251) );
  NAND2X0 U1751 ( .IN1(n256), .IN2(n12), .QN(n254) );
  NAND2X0 U1752 ( .IN1(n259), .IN2(n12), .QN(n257) );
  NAND2X0 U1761 ( .IN1(n262), .IN2(n12), .QN(n260) );
  NAND2X0 U1762 ( .IN1(n265), .IN2(n12), .QN(n263) );
  NAND2X0 U1771 ( .IN1(n268), .IN2(n9), .QN(n266) );
  NAND2X0 U1772 ( .IN1(n271), .IN2(n9), .QN(n269) );
  NAND2X0 U1781 ( .IN1(n274), .IN2(n9), .QN(n272) );
  NAND2X0 U1782 ( .IN1(n277), .IN2(n9), .QN(n275) );
  NAND2X0 U1791 ( .IN1(n280), .IN2(n9), .QN(n278) );
  NAND2X0 U1792 ( .IN1(n283), .IN2(n9), .QN(n281) );
  NAND2X0 U1801 ( .IN1(n286), .IN2(n9), .QN(n284) );
  NAND2X0 U1802 ( .IN1(n289), .IN2(n9), .QN(n287) );
  NAND2X0 U1811 ( .IN1(n292), .IN2(n9), .QN(n290) );
  NAND2X0 U1812 ( .IN1(n295), .IN2(n9), .QN(n293) );
  NAND2X0 U1821 ( .IN1(n298), .IN2(n9), .QN(n296) );
  NAND2X0 U1822 ( .IN1(n301), .IN2(n9), .QN(n299) );
  NAND2X0 U1831 ( .IN1(n304), .IN2(n6), .QN(n302) );
  NAND2X0 U1832 ( .IN1(n307), .IN2(n6), .QN(n305) );
  NAND2X0 U1841 ( .IN1(n310), .IN2(n6), .QN(n308) );
  NAND2X0 U1842 ( .IN1(n313), .IN2(n6), .QN(n311) );
  NAND2X0 U1851 ( .IN1(n316), .IN2(n6), .QN(n314) );
  NAND2X0 U1852 ( .IN1(n319), .IN2(n6), .QN(n317) );
  NAND2X0 U1861 ( .IN1(n322), .IN2(n6), .QN(n320) );
  NAND2X0 U1862 ( .IN1(n325), .IN2(n6), .QN(n323) );
  NAND2X0 U1871 ( .IN1(n328), .IN2(n6), .QN(n326) );
  NAND2X0 U1872 ( .IN1(n331), .IN2(n6), .QN(n329) );
  NAND2X0 U1881 ( .IN1(n334), .IN2(n6), .QN(n332) );
  NAND2X0 U1882 ( .IN1(n337), .IN2(n6), .QN(n335) );
  NAND2X0 U1891 ( .IN1(n340), .IN2(n2), .QN(n338) );
  NAND2X0 U1892 ( .IN1(n343), .IN2(n2), .QN(n341) );
  NAND2X0 U1901 ( .IN1(n346), .IN2(n2), .QN(n344) );
  NAND2X0 U1902 ( .IN1(n349), .IN2(n2), .QN(n347) );
  NAND2X0 U1911 ( .IN1(n352), .IN2(n2), .QN(n350) );
  NAND2X0 U1912 ( .IN1(n355), .IN2(n2), .QN(n353) );
  NAND2X0 U1921 ( .IN1(n358), .IN2(n2), .QN(n356) );
  NAND2X0 U1922 ( .IN1(n361), .IN2(n2), .QN(n359) );
  NAND2X0 U1931 ( .IN1(n364), .IN2(n2), .QN(n362) );
  NAND2X0 U1932 ( .IN1(n367), .IN2(n2), .QN(n365) );
  NAND2X0 U1941 ( .IN1(n370), .IN2(n2), .QN(n368) );
  NAND2X0 U1942 ( .IN1(n373), .IN2(n2), .QN(n371) );
  NAND2X0 U1951 ( .IN1(n376), .IN2(n9), .QN(n374) );
  NAND2X0 U1952 ( .IN1(n379), .IN2(n6), .QN(n377) );
  NAND2X0 U1961 ( .IN1(n382), .IN2(n2), .QN(n380) );
  NAND2X0 U1962 ( .IN1(n385), .IN2(n9), .QN(n383) );
  NAND2X0 U1971 ( .IN1(n388), .IN2(n6), .QN(n386) );
  NAND2X0 U1972 ( .IN1(n391), .IN2(n2), .QN(n389) );
  NAND2X0 U1981 ( .IN1(n394), .IN2(n30), .QN(n392) );
  NAND2X0 U1982 ( .IN1(n397), .IN2(n2), .QN(n395) );
  NAND2X0 U1991 ( .IN1(n400), .IN2(n27), .QN(n398) );
  NAND2X0 U1992 ( .IN1(n403), .IN2(n2), .QN(n401) );
  NAND2X0 U2001 ( .IN1(n406), .IN2(n4), .QN(n404) );
  NAND2X0 U2002 ( .IN1(n409), .IN2(n30), .QN(n407) );
  NAND2X0 U2011 ( .IN1(n412), .IN2(n18), .QN(n410) );
  NAND2X0 U2012 ( .IN1(n415), .IN2(n24), .QN(n413) );
  NAND2X0 U2021 ( .IN1(n418), .IN2(n9), .QN(n416) );
  NAND2X0 U2022 ( .IN1(n421), .IN2(n2), .QN(n419) );
  NAND2X0 U2031 ( .IN1(n424), .IN2(n6), .QN(n422) );
  NAND2X0 U2032 ( .IN1(n427), .IN2(n6), .QN(n425) );
  NAND2X0 U2041 ( .IN1(n430), .IN2(n21), .QN(n428) );
  NAND2X0 U2042 ( .IN1(n433), .IN2(n4), .QN(n431) );
  NAND2X0 U2051 ( .IN1(n436), .IN2(n30), .QN(n434) );
  NAND2X0 U2052 ( .IN1(n439), .IN2(n12), .QN(n437) );
  NAND2X0 U2061 ( .IN1(n442), .IN2(n6), .QN(n440) );
  NAND2X0 U2062 ( .IN1(n445), .IN2(n2), .QN(n443) );
  NAND2X0 U2071 ( .IN1(n448), .IN2(n9), .QN(n446) );
  NAND2X0 U2072 ( .IN1(n451), .IN2(n6), .QN(n449) );
  NAND2X0 U2081 ( .IN1(n454), .IN2(n4), .QN(n452) );
  NAND2X0 U2082 ( .IN1(n457), .IN2(n4), .QN(n455) );
  NAND2X0 U2091 ( .IN1(n460), .IN2(n4), .QN(n458) );
  NAND2X0 U2092 ( .IN1(n463), .IN2(n4), .QN(n461) );
  NAND2X0 U2101 ( .IN1(n466), .IN2(n4), .QN(n464) );
  NAND2X0 U2102 ( .IN1(n469), .IN2(n4), .QN(n467) );
  NAND2X0 U2111 ( .IN1(n472), .IN2(n4), .QN(n470) );
  NAND2X0 U2112 ( .IN1(n475), .IN2(n4), .QN(n473) );
  NAND2X0 U2121 ( .IN1(n478), .IN2(n4), .QN(n476) );
  NAND2X0 U2122 ( .IN1(n481), .IN2(n4), .QN(n479) );
  NAND2X0 U2131 ( .IN1(n484), .IN2(n18), .QN(n482) );
  NAND2X0 U2132 ( .IN1(n487), .IN2(n15), .QN(n485) );
  NAND2X0 U2141 ( .IN1(n490), .IN2(n12), .QN(n488) );
  NAND2X0 U2142 ( .IN1(n493), .IN2(n9), .QN(n491) );
  NAND2X0 U2151 ( .IN1(n496), .IN2(n4), .QN(n494) );
  NAND2X0 U2152 ( .IN1(n499), .IN2(n4), .QN(n497) );
  NAND2X0 U2161 ( .IN1(n502), .IN2(n4), .QN(n500) );
  NAND2X0 U2162 ( .IN1(n505), .IN2(n4), .QN(n503) );
  NAND2X0 U2171 ( .IN1(n508), .IN2(n4), .QN(n506) );
  NAND2X0 U2172 ( .IN1(n511), .IN2(n4), .QN(n509) );
  NAND2X0 U2181 ( .IN1(n514), .IN2(n4), .QN(n512) );
  NAND2X0 U2182 ( .IN1(n517), .IN2(n4), .QN(n515) );
  NAND2X0 U2191 ( .IN1(n520), .IN2(n27), .QN(n518) );
  NAND2X0 U2192 ( .IN1(n523), .IN2(n24), .QN(n521) );
  NAND2X0 U2201 ( .IN1(n526), .IN2(n21), .QN(n524) );
  NAND2X0 U2202 ( .IN1(n529), .IN2(n18), .QN(n527) );
  NAND2X0 U2211 ( .IN1(n532), .IN2(n15), .QN(n530) );
  NAND2X0 U2212 ( .IN1(n535), .IN2(n12), .QN(n533) );
  NAND2X0 U2221 ( .IN1(n538), .IN2(n30), .QN(n536) );
  NAND2X0 U2222 ( .IN1(n541), .IN2(n27), .QN(n539) );
  NAND2X0 U2231 ( .IN1(n544), .IN2(n24), .QN(n542) );
  NAND2X0 U2232 ( .IN1(n547), .IN2(n21), .QN(n545) );
  NAND2X0 U2241 ( .IN1(n550), .IN2(n18), .QN(n548) );
  NAND2X0 U2242 ( .IN1(n553), .IN2(n15), .QN(n551) );
  NAND2X0 U2251 ( .IN1(n556), .IN2(n24), .QN(n554) );
  NAND2X0 U2252 ( .IN1(n559), .IN2(n21), .QN(n557) );
  NAND2X0 U2261 ( .IN1(n562), .IN2(n18), .QN(n560) );
  NAND2X0 U2262 ( .IN1(n565), .IN2(n15), .QN(n563) );
  NAND2X0 U2271 ( .IN1(n568), .IN2(n12), .QN(n566) );
  NAND2X0 U2272 ( .IN1(n571), .IN2(n9), .QN(n569) );
  NAND2X0 U2281 ( .IN1(n574), .IN2(n4), .QN(n572) );
  NAND2X0 U2282 ( .IN1(n577), .IN2(n4), .QN(n575) );
  NAND2X0 U2291 ( .IN1(n580), .IN2(n4), .QN(n578) );
  NAND2X0 U2292 ( .IN1(n583), .IN2(n4), .QN(n581) );
  NAND2X0 U2301 ( .IN1(n586), .IN2(n4), .QN(n584) );
  NAND2X0 U2302 ( .IN1(n589), .IN2(n4), .QN(n587) );
  NAND2X0 U2311 ( .IN1(n592), .IN2(n30), .QN(n590) );
  NAND2X0 U2312 ( .IN1(n595), .IN2(n27), .QN(n593) );
  NAND2X0 U2321 ( .IN1(n598), .IN2(n24), .QN(n596) );
  NAND2X0 U2322 ( .IN1(n601), .IN2(n21), .QN(n599) );
  NAND2X0 U2331 ( .IN1(n604), .IN2(n18), .QN(n602) );
  NAND2X0 U2332 ( .IN1(n607), .IN2(n15), .QN(n605) );
  NAND2X0 U2341 ( .IN1(n610), .IN2(n12), .QN(n608) );
  NAND2X0 U2342 ( .IN1(n613), .IN2(n9), .QN(n611) );
  NAND2X0 U2351 ( .IN1(n616), .IN2(n4), .QN(n614) );
  NAND2X0 U2352 ( .IN1(n619), .IN2(n4), .QN(n617) );
  NAND2X0 U2361 ( .IN1(n622), .IN2(n4), .QN(n620) );
  NAND2X0 U2362 ( .IN1(n625), .IN2(n4), .QN(n623) );
  NAND2X0 U2371 ( .IN1(n628), .IN2(n2), .QN(n626) );
  NAND2X0 U2372 ( .IN1(n631), .IN2(n2), .QN(n629) );
  NAND2X0 U2381 ( .IN1(n634), .IN2(n30), .QN(n632) );
  NAND2X0 U2382 ( .IN1(n637), .IN2(n27), .QN(n635) );
  NAND2X0 U2391 ( .IN1(n640), .IN2(n24), .QN(n638) );
  NAND2X0 U2392 ( .IN1(n643), .IN2(n21), .QN(n641) );
  NAND2X0 U2401 ( .IN1(n646), .IN2(n18), .QN(n644) );
  NAND2X0 U2402 ( .IN1(n649), .IN2(n15), .QN(n647) );
  NAND2X0 U2411 ( .IN1(n652), .IN2(n12), .QN(n650) );
  NAND2X0 U2412 ( .IN1(n655), .IN2(n9), .QN(n653) );
  NAND2X0 U2421 ( .IN1(n658), .IN2(n4), .QN(n656) );
  NAND2X0 U2422 ( .IN1(n661), .IN2(n4), .QN(n659) );
  NAND2X0 U2431 ( .IN1(n664), .IN2(n24), .QN(n662) );
  NAND2X0 U2432 ( .IN1(n667), .IN2(n6), .QN(n665) );
  NAND2X0 U2441 ( .IN1(n670), .IN2(n2), .QN(n668) );
  NAND2X0 U2442 ( .IN1(n673), .IN2(n27), .QN(n671) );
  NAND2X0 U2451 ( .IN1(n676), .IN2(n30), .QN(n674) );
  NAND2X0 U2452 ( .IN1(n679), .IN2(n27), .QN(n677) );
  NAND2X0 U2461 ( .IN1(n682), .IN2(n24), .QN(n680) );
  NAND2X0 U2462 ( .IN1(n685), .IN2(n21), .QN(n683) );
  NAND2X0 U2471 ( .IN1(n688), .IN2(n18), .QN(n686) );
  NAND2X0 U2472 ( .IN1(n691), .IN2(n15), .QN(n689) );
  NAND2X0 U2481 ( .IN1(n694), .IN2(n12), .QN(n692) );
  NAND2X0 U2482 ( .IN1(n697), .IN2(n9), .QN(n695) );
  NAND2X0 U2491 ( .IN1(n700), .IN2(n4), .QN(n698) );
  NAND2X0 U2492 ( .IN1(n703), .IN2(n4), .QN(n701) );
  NAND2X0 U2501 ( .IN1(n706), .IN2(n4), .QN(n704) );
  NAND2X0 U2502 ( .IN1(n709), .IN2(n4), .QN(n707) );
  NAND2X0 U2511 ( .IN1(n712), .IN2(n4), .QN(n710) );
  NAND2X0 U2512 ( .IN1(n715), .IN2(n4), .QN(n713) );
  NAND2X0 U2521 ( .IN1(n718), .IN2(n4), .QN(n716) );
  NAND2X0 U2522 ( .IN1(n721), .IN2(n4), .QN(n719) );
  NAND2X0 U2531 ( .IN1(n724), .IN2(n4), .QN(n722) );
  NAND2X0 U2532 ( .IN1(n727), .IN2(n4), .QN(n725) );
  NAND2X0 U2541 ( .IN1(n730), .IN2(n4), .QN(n728) );
  NAND2X0 U2542 ( .IN1(n733), .IN2(n4), .QN(n731) );
  NAND2X0 U2551 ( .IN1(n736), .IN2(n27), .QN(n734) );
  NAND2X0 U2552 ( .IN1(n739), .IN2(n6), .QN(n737) );
  NAND2X0 U2561 ( .IN1(n742), .IN2(n6), .QN(n740) );
  NAND2X0 U2562 ( .IN1(n745), .IN2(n30), .QN(n743) );
  NAND2X0 U2563 ( .IN1(n748), .IN2(n4), .QN(n746) );
  NAND2X0 U2566 ( .IN1(n751), .IN2(n30), .QN(n749) );
  NAND2X0 U2603 ( .IN1(n754), .IN2(n27), .QN(n752) );
  NAND2X0 U2640 ( .IN1(n757), .IN2(n24), .QN(n755) );
  NAND2X0 U2677 ( .IN1(n760), .IN2(n21), .QN(n758) );
  NAND2X0 U2716 ( .IN1(n763), .IN2(n18), .QN(n761) );
  NAND2X0 U2753 ( .IN1(n766), .IN2(n15), .QN(n764) );
  NAND2X0 U2790 ( .IN1(n769), .IN2(n12), .QN(n767) );
  NAND2X0 U2827 ( .IN1(n7), .IN2(n21), .QN(n5) );
  NAND2X0 U2866 ( .IN1(n10), .IN2(n15), .QN(n8) );
  NAND2X0 U2903 ( .IN1(n13), .IN2(n12), .QN(n11) );
  INVX0 U2940 ( .IN(n4), .QN(n33) );
  INVX0 U2977 ( .IN(n771), .QN(n4174) );
  AND2X1 U3016 ( .IN1(n1843), .IN2(n1862), .Q(n3) );
  NOR2X0 U3053 ( .IN1(n4175), .IN2(R), .QN(n4) );
  AND2X1 U3090 ( .IN1(n1964), .IN2(n1943), .Q(n1862) );
  AND2X1 U3127 ( .IN1(n1962), .IN2(n1921), .Q(n1843) );
  NAND2X0 U3166 ( .IN1(R), .IN2(n4175), .QN(n771) );
  AND2X1 U3203 ( .IN1(n1850), .IN2(n1833), .Q(n355) );
  AND2X1 U3240 ( .IN1(n1853), .IN2(n1833), .Q(n307) );
  AND2X1 U3277 ( .IN1(n1850), .IN2(n1838), .Q(n379) );
  AND2X1 U3316 ( .IN1(n1853), .IN2(n1838), .Q(n331) );
  AND2X1 U3353 ( .IN1(n1829), .IN2(n1833), .Q(n259) );
  AND2X1 U3390 ( .IN1(n1842), .IN2(n1833), .Q(n211) );
  AND2X1 U3427 ( .IN1(n1829), .IN2(n1838), .Q(n283) );
  AND2X1 U3466 ( .IN1(n1842), .IN2(n1838), .Q(n235) );
  AND2X1 U3503 ( .IN1(n1861), .IN2(n1831), .Q(n106) );
  AND2X1 U3540 ( .IN1(n1840), .IN2(n1837), .Q(n190) );
  AND2X1 U3577 ( .IN1(n1840), .IN2(n1832), .Q(n166) );
  AND2X1 U3616 ( .IN1(n1861), .IN2(n1837), .Q(n142) );
  AND2X1 U3620 ( .IN1(n1860), .IN2(n1832), .Q(n70) );
  AND2X1 U3621 ( .IN1(n1860), .IN2(n1837), .Q(n94) );
  AND2X1 U3622 ( .IN1(n1838), .IN2(n1862), .Q(n43) );
  AND2X1 U3623 ( .IN1(n1866), .IN2(n1862), .Q(n13) );
  AND2X1 U3626 ( .IN1(n1915), .IN2(n1833), .Q(n547) );
  AND2X1 U3627 ( .IN1(n1918), .IN2(n1833), .Q(n499) );
  AND2X1 U3628 ( .IN1(n1915), .IN2(n1838), .Q(n571) );
  AND2X1 U3629 ( .IN1(n1918), .IN2(n1838), .Q(n523) );
  AND2X1 U3632 ( .IN1(n1873), .IN2(n1833), .Q(n739) );
  AND2X1 U3633 ( .IN1(n1898), .IN2(n1833), .Q(n691) );
  AND2X1 U3634 ( .IN1(n1873), .IN2(n1838), .Q(n763) );
  AND2X1 U3635 ( .IN1(n1898), .IN2(n1838), .Q(n715) );
  AND2X1 U3638 ( .IN1(n1886), .IN2(n1833), .Q(n643) );
  AND2X1 U3639 ( .IN1(n1889), .IN2(n1833), .Q(n595) );
  AND2X1 U3640 ( .IN1(n1886), .IN2(n1838), .Q(n667) );
  AND2X1 U3641 ( .IN1(n1889), .IN2(n1838), .Q(n619) );
  AND2X1 U3645 ( .IN1(n1905), .IN2(n1833), .Q(n451) );
  AND2X1 U3646 ( .IN1(n1908), .IN2(n1833), .Q(n403) );
  AND2X1 U3647 ( .IN1(n1905), .IN2(n1838), .Q(n475) );
  AND2X1 U3648 ( .IN1(n1908), .IN2(n1838), .Q(n427) );
  AND2X1 U3651 ( .IN1(n1840), .IN2(n1866), .Q(n157) );
  AND2X1 U3652 ( .IN1(n1840), .IN2(n1939), .Q(n181) );
  AND2X1 U3653 ( .IN1(n1861), .IN2(n1866), .Q(n109) );
  AND2X1 U3654 ( .IN1(n1861), .IN2(n1939), .Q(n133) );
  AND2X1 U3657 ( .IN1(n1850), .IN2(n1866), .Q(n349) );
  AND2X1 U3658 ( .IN1(n1850), .IN2(n1939), .Q(n373) );
  AND2X1 U3659 ( .IN1(n1853), .IN2(n1866), .Q(n301) );
  AND2X1 U3660 ( .IN1(n1853), .IN2(n1939), .Q(n325) );
  AND2X1 U3663 ( .IN1(n1829), .IN2(n1866), .Q(n253) );
  AND2X1 U3664 ( .IN1(n1829), .IN2(n1939), .Q(n277) );
  AND2X1 U3665 ( .IN1(n1842), .IN2(n1866), .Q(n205) );
  AND2X1 U3666 ( .IN1(n1842), .IN2(n1939), .Q(n229) );
  AND2X1 U3670 ( .IN1(n1860), .IN2(n1866), .Q(n61) );
  AND2X1 U3671 ( .IN1(n1860), .IN2(n1939), .Q(n85) );
  AND2X1 U3672 ( .IN1(n1833), .IN2(n1862), .Q(n19) );
  AND2X1 U3673 ( .IN1(n1939), .IN2(n1862), .Q(n37) );
  AND2X1 U3676 ( .IN1(n1915), .IN2(n1866), .Q(n541) );
  AND2X1 U3677 ( .IN1(n1915), .IN2(n1939), .Q(n565) );
  AND2X1 U3678 ( .IN1(n1918), .IN2(n1866), .Q(n493) );
  AND2X1 U3679 ( .IN1(n1918), .IN2(n1939), .Q(n517) );
  AND2X1 U3682 ( .IN1(n1873), .IN2(n1866), .Q(n733) );
  AND2X1 U3683 ( .IN1(n1873), .IN2(n1939), .Q(n757) );
  AND2X1 U3684 ( .IN1(n1898), .IN2(n1866), .Q(n685) );
  AND2X1 U3685 ( .IN1(n1898), .IN2(n1939), .Q(n709) );
  AND2X1 U3688 ( .IN1(n1886), .IN2(n1866), .Q(n637) );
  AND2X1 U3689 ( .IN1(n1886), .IN2(n1939), .Q(n661) );
  AND2X1 U3690 ( .IN1(n1889), .IN2(n1866), .Q(n589) );
  AND2X1 U3691 ( .IN1(n1889), .IN2(n1939), .Q(n613) );
  AND2X1 U3695 ( .IN1(n1905), .IN2(n1866), .Q(n445) );
  AND2X1 U3696 ( .IN1(n1905), .IN2(n1939), .Q(n469) );
  AND2X1 U3697 ( .IN1(n1908), .IN2(n1866), .Q(n397) );
  AND2X1 U3698 ( .IN1(n1908), .IN2(n1939), .Q(n421) );
  AND2X1 U3701 ( .IN1(n1850), .IN2(n1831), .Q(n346) );
  AND2X1 U3702 ( .IN1(n1853), .IN2(n1831), .Q(n298) );
  AND2X1 U3703 ( .IN1(n1850), .IN2(n1836), .Q(n370) );
  AND2X1 U3704 ( .IN1(n1853), .IN2(n1836), .Q(n322) );
  AND2X1 U3707 ( .IN1(n1829), .IN2(n1831), .Q(n250) );
  AND2X1 U3708 ( .IN1(n1842), .IN2(n1843), .Q(n196) );
  AND2X1 U3709 ( .IN1(n1829), .IN2(n1836), .Q(n274) );
  AND2X1 U3710 ( .IN1(n1842), .IN2(n1836), .Q(n226) );
  AND2X1 U3713 ( .IN1(n1861), .IN2(n1830), .Q(n103) );
  AND2X1 U3714 ( .IN1(n1840), .IN2(n1833), .Q(n163) );
  AND2X1 U3715 ( .IN1(n1873), .IN2(n1841), .Q(n769) );
  AND2X1 U3716 ( .IN1(n1861), .IN2(n1833), .Q(n115) );
  AND2X1 U3717 ( .IN1(n1861), .IN2(n1838), .Q(n139) );
  AND2X1 U3721 ( .IN1(n1860), .IN2(n1833), .Q(n67) );
  AND2X1 U3722 ( .IN1(n1836), .IN2(n1862), .Q(n34) );
  AND2X1 U3723 ( .IN1(n1860), .IN2(n1838), .Q(n91) );
  AND2X1 U3724 ( .IN1(n1915), .IN2(n1831), .Q(n538) );
  AND2X1 U3727 ( .IN1(n1918), .IN2(n1831), .Q(n490) );
  AND2X1 U3728 ( .IN1(n1915), .IN2(n1836), .Q(n562) );
  AND2X1 U3729 ( .IN1(n1918), .IN2(n1836), .Q(n514) );
  AND2X1 U3730 ( .IN1(n1873), .IN2(n1831), .Q(n730) );
  AND2X1 U3733 ( .IN1(n1898), .IN2(n1831), .Q(n682) );
  AND2X1 U3734 ( .IN1(n1873), .IN2(n1836), .Q(n754) );
  AND2X1 U3735 ( .IN1(n1898), .IN2(n1836), .Q(n706) );
  AND2X1 U3736 ( .IN1(n1886), .IN2(n1831), .Q(n634) );
  AND2X1 U3739 ( .IN1(n1889), .IN2(n1831), .Q(n586) );
  AND2X1 U3740 ( .IN1(n1886), .IN2(n1836), .Q(n658) );
  AND2X1 U3741 ( .IN1(n1889), .IN2(n1836), .Q(n610) );
  AND2X1 U3742 ( .IN1(n1905), .IN2(n1831), .Q(n442) );
  AND2X1 U3746 ( .IN1(n1908), .IN2(n1831), .Q(n394) );
  AND2X1 U3747 ( .IN1(n1905), .IN2(n1836), .Q(n466) );
  AND2X1 U3748 ( .IN1(n1908), .IN2(n1836), .Q(n418) );
  AND2X1 U3749 ( .IN1(n1840), .IN2(n1843), .Q(n148) );
  AND2X1 U3752 ( .IN1(n1840), .IN2(n1937), .Q(n172) );
  AND2X1 U3753 ( .IN1(n1861), .IN2(n1843), .Q(n100) );
  AND2X1 U3754 ( .IN1(n1861), .IN2(n1937), .Q(n124) );
  AND2X1 U3755 ( .IN1(n1850), .IN2(n1843), .Q(n340) );
  AND2X1 U3758 ( .IN1(n1850), .IN2(n1937), .Q(n364) );
  AND2X1 U3759 ( .IN1(n1853), .IN2(n1843), .Q(n292) );
  AND2X1 U3760 ( .IN1(n1853), .IN2(n1937), .Q(n316) );
  AND2X1 U3761 ( .IN1(n1829), .IN2(n1843), .Q(n244) );
  AND2X1 U3764 ( .IN1(n1829), .IN2(n1937), .Q(n268) );
  AND2X1 U3765 ( .IN1(n1842), .IN2(n1831), .Q(n202) );
  AND2X1 U3766 ( .IN1(n1842), .IN2(n1937), .Q(n220) );
  AND2X1 U3767 ( .IN1(n1860), .IN2(n1831), .Q(n58) );
  AND2X1 U3771 ( .IN1(n1860), .IN2(n1937), .Q(n76) );
  AND2X1 U3772 ( .IN1(n1831), .IN2(n1862), .Q(n10) );
  AND2X1 U3773 ( .IN1(n1937), .IN2(n1862), .Q(n28) );
  AND2X1 U3774 ( .IN1(n1915), .IN2(n1843), .Q(n532) );
  AND2X1 U3777 ( .IN1(n1915), .IN2(n1937), .Q(n556) );
  AND2X1 U3778 ( .IN1(n1918), .IN2(n1843), .Q(n484) );
  AND2X1 U3779 ( .IN1(n1918), .IN2(n1937), .Q(n508) );
  AND2X1 U3780 ( .IN1(n1873), .IN2(n1843), .Q(n724) );
  AND2X1 U3783 ( .IN1(n1873), .IN2(n1937), .Q(n748) );
  AND2X1 U3784 ( .IN1(n1898), .IN2(n1843), .Q(n676) );
  AND2X1 U3785 ( .IN1(n1898), .IN2(n1937), .Q(n700) );
  AND2X1 U3786 ( .IN1(n1886), .IN2(n1843), .Q(n628) );
  AND2X1 U3789 ( .IN1(n1886), .IN2(n1937), .Q(n652) );
  AND2X1 U3790 ( .IN1(n1889), .IN2(n1843), .Q(n580) );
  AND2X1 U3791 ( .IN1(n1889), .IN2(n1937), .Q(n604) );
  AND2X1 U3792 ( .IN1(n1905), .IN2(n1843), .Q(n436) );
  AND2X1 U3796 ( .IN1(n1905), .IN2(n1937), .Q(n460) );
  AND2X1 U3797 ( .IN1(n1908), .IN2(n1843), .Q(n388) );
  AND2X1 U3798 ( .IN1(n1908), .IN2(n1937), .Q(n412) );
  AND2X1 U3799 ( .IN1(n1850), .IN2(n1830), .Q(n343) );
  AND2X1 U3802 ( .IN1(n1853), .IN2(n1830), .Q(n295) );
  AND2X1 U3803 ( .IN1(n1850), .IN2(n1835), .Q(n367) );
  AND2X1 U3804 ( .IN1(n1853), .IN2(n1835), .Q(n319) );
  AND2X1 U3805 ( .IN1(n1829), .IN2(n1830), .Q(n247) );
  AND2X1 U3808 ( .IN1(n1840), .IN2(n1841), .Q(n193) );
  AND2X1 U3809 ( .IN1(n1829), .IN2(n1835), .Q(n271) );
  AND2X1 U3810 ( .IN1(n1842), .IN2(n1835), .Q(n223) );
  AND2X1 U3811 ( .IN1(n1861), .IN2(n1832), .Q(n118) );
  AND2X1 U3814 ( .IN1(n1840), .IN2(n1836), .Q(n178) );
  AND2X1 U3815 ( .IN1(n1840), .IN2(n1831), .Q(n154) );
  AND2X1 U3816 ( .IN1(n1861), .IN2(n1836), .Q(n130) );
  AND2X1 U3817 ( .IN1(n1860), .IN2(n1843), .Q(n52) );
  AND2X1 U3818 ( .IN1(n1860), .IN2(n1836), .Q(n82) );
  AND2X1 U3819 ( .IN1(n1835), .IN2(n1862), .Q(n31) );
  AND2X1 U3820 ( .IN1(n1915), .IN2(n1830), .Q(n535) );
  AND2X1 U3821 ( .IN1(n1918), .IN2(n1830), .Q(n487) );
  AND2X1 U3822 ( .IN1(n1915), .IN2(n1835), .Q(n559) );
  AND2X1 U3826 ( .IN1(n1918), .IN2(n1835), .Q(n511) );
  AND2X1 U3827 ( .IN1(n1873), .IN2(n1830), .Q(n727) );
  AND2X1 U3828 ( .IN1(n1898), .IN2(n1830), .Q(n679) );
  AND2X1 U3829 ( .IN1(n1873), .IN2(n1835), .Q(n751) );
  AND2X1 U3832 ( .IN1(n1898), .IN2(n1835), .Q(n703) );
  AND2X1 U3833 ( .IN1(n1886), .IN2(n1830), .Q(n631) );
  AND2X1 U3834 ( .IN1(n1889), .IN2(n1830), .Q(n583) );
  AND2X1 U3835 ( .IN1(n1886), .IN2(n1835), .Q(n655) );
  AND2X1 U3838 ( .IN1(n1889), .IN2(n1835), .Q(n607) );
  AND2X1 U3839 ( .IN1(n1905), .IN2(n1830), .Q(n439) );
  AND2X1 U3840 ( .IN1(n1908), .IN2(n1830), .Q(n391) );
  AND2X1 U3841 ( .IN1(n1905), .IN2(n1835), .Q(n463) );
  AND2X1 U3844 ( .IN1(n1908), .IN2(n1835), .Q(n415) );
  AND2X1 U3845 ( .IN1(n1861), .IN2(n1841), .Q(n145) );
  AND2X1 U3846 ( .IN1(n1840), .IN2(n1936), .Q(n169) );
  AND2X1 U3847 ( .IN1(n1860), .IN2(n1841), .Q(n97) );
  AND2X1 U3848 ( .IN1(n1861), .IN2(n1936), .Q(n121) );
  AND2X1 U3852 ( .IN1(n1853), .IN2(n1841), .Q(n337) );
  AND2X1 U3853 ( .IN1(n1850), .IN2(n1936), .Q(n361) );
  AND2X1 U3854 ( .IN1(n1829), .IN2(n1841), .Q(n289) );
  AND2X1 U3855 ( .IN1(n1853), .IN2(n1936), .Q(n313) );
  AND2X1 U3858 ( .IN1(n1842), .IN2(n1841), .Q(n241) );
  AND2X1 U3859 ( .IN1(n1829), .IN2(n1936), .Q(n265) );
  AND2X1 U3860 ( .IN1(n1842), .IN2(n1830), .Q(n199) );
  AND2X1 U3861 ( .IN1(n1842), .IN2(n1936), .Q(n217) );
  AND2X1 U3864 ( .IN1(n1860), .IN2(n1830), .Q(n55) );
  AND2X1 U3865 ( .IN1(n1860), .IN2(n1936), .Q(n73) );
  AND2X1 U3866 ( .IN1(n1830), .IN2(n1862), .Q(n7) );
  AND2X1 U3867 ( .IN1(n1936), .IN2(n1862), .Q(n25) );
  AND2X1 U3868 ( .IN1(n1918), .IN2(n1841), .Q(n529) );
  AND2X1 U3871 ( .IN1(n1915), .IN2(n1936), .Q(n553) );
  AND2X1 U3872 ( .IN1(n1905), .IN2(n1841), .Q(n481) );
  AND2X1 U3873 ( .IN1(n1918), .IN2(n1936), .Q(n505) );
  AND2X1 U3874 ( .IN1(n1898), .IN2(n1841), .Q(n721) );
  AND2X1 U3875 ( .IN1(n1873), .IN2(n1936), .Q(n745) );
  AND2X1 U3879 ( .IN1(n1886), .IN2(n1841), .Q(n673) );
  AND2X1 U3880 ( .IN1(n1898), .IN2(n1936), .Q(n697) );
  AND2X1 U3881 ( .IN1(n1889), .IN2(n1841), .Q(n625) );
  AND2X1 U3882 ( .IN1(n1886), .IN2(n1936), .Q(n649) );
  AND2X1 U3885 ( .IN1(n1915), .IN2(n1841), .Q(n577) );
  AND2X1 U3886 ( .IN1(n1889), .IN2(n1936), .Q(n601) );
  AND2X1 U3887 ( .IN1(n1908), .IN2(n1841), .Q(n433) );
  AND2X1 U3888 ( .IN1(n1905), .IN2(n1936), .Q(n457) );
  AND2X1 U3891 ( .IN1(n1850), .IN2(n1841), .Q(n385) );
  AND2X1 U3892 ( .IN1(n1908), .IN2(n1936), .Q(n409) );
  AND2X1 U3893 ( .IN1(n1850), .IN2(n1832), .Q(n358) );
  AND2X1 U3894 ( .IN1(n1853), .IN2(n1832), .Q(n310) );
  AND2X1 U3895 ( .IN1(n1850), .IN2(n1837), .Q(n382) );
  AND2X1 U3896 ( .IN1(n1853), .IN2(n1837), .Q(n334) );
  AND2X1 U3897 ( .IN1(n1829), .IN2(n1832), .Q(n262) );
  AND2X1 U3898 ( .IN1(n1842), .IN2(n1832), .Q(n214) );
  AND2X1 U3901 ( .IN1(n1829), .IN2(n1837), .Q(n286) );
  AND2X1 U3902 ( .IN1(n1842), .IN2(n1837), .Q(n238) );
  AND2X1 U3903 ( .IN1(n1840), .IN2(n1838), .Q(n187) );
  AND2X1 U3904 ( .IN1(n1840), .IN2(n1835), .Q(n175) );
  AND2X1 U3905 ( .IN1(n1840), .IN2(n1830), .Q(n151) );
  AND2X1 U3909 ( .IN1(n1861), .IN2(n1835), .Q(n127) );
  AND2X1 U3910 ( .IN1(n1841), .IN2(n1862), .Q(n49) );
  AND2X1 U3911 ( .IN1(n1860), .IN2(n1835), .Q(n79) );
  AND2X1 U3912 ( .IN1(n1837), .IN2(n1862), .Q(n46) );
  AND2X1 U3915 ( .IN1(n1865), .IN2(n1862), .Q(n16) );
  AND2X1 U3916 ( .IN1(n1915), .IN2(n1832), .Q(n550) );
  AND2X1 U3917 ( .IN1(n1918), .IN2(n1832), .Q(n502) );
  AND2X1 U3918 ( .IN1(n1915), .IN2(n1837), .Q(n574) );
  AND2X1 U3919 ( .IN1(n1918), .IN2(n1837), .Q(n526) );
  AND2X1 U3922 ( .IN1(n1873), .IN2(n1832), .Q(n742) );
  AND2X1 U3923 ( .IN1(n1898), .IN2(n1832), .Q(n694) );
  AND2X1 U3924 ( .IN1(n1873), .IN2(n1837), .Q(n766) );
  AND2X1 U3925 ( .IN1(n1898), .IN2(n1837), .Q(n718) );
  AND2X1 U3926 ( .IN1(n1886), .IN2(n1832), .Q(n646) );
  AND2X1 U3929 ( .IN1(n1889), .IN2(n1832), .Q(n598) );
  AND2X1 U3930 ( .IN1(n1886), .IN2(n1837), .Q(n670) );
  AND2X1 U3931 ( .IN1(n1889), .IN2(n1837), .Q(n622) );
  AND2X1 U3932 ( .IN1(n1905), .IN2(n1832), .Q(n454) );
  AND2X1 U3933 ( .IN1(n1908), .IN2(n1832), .Q(n406) );
  AND2X1 U3934 ( .IN1(n1905), .IN2(n1837), .Q(n478) );
  AND2X1 U3935 ( .IN1(n1908), .IN2(n1837), .Q(n430) );
  AND2X1 U3939 ( .IN1(n1840), .IN2(n1865), .Q(n160) );
  AND2X1 U3940 ( .IN1(n1840), .IN2(n1938), .Q(n184) );
  AND2X1 U3941 ( .IN1(n1861), .IN2(n1865), .Q(n112) );
  AND2X1 U3942 ( .IN1(n1861), .IN2(n1938), .Q(n136) );
  AND2X1 U3945 ( .IN1(n1850), .IN2(n1865), .Q(n352) );
  AND2X1 U3946 ( .IN1(n1850), .IN2(n1938), .Q(n376) );
  AND2X1 U3947 ( .IN1(n1853), .IN2(n1865), .Q(n304) );
  AND2X1 U3948 ( .IN1(n1853), .IN2(n1938), .Q(n328) );
  AND2X1 U3951 ( .IN1(n1829), .IN2(n1865), .Q(n256) );
  AND2X1 U3952 ( .IN1(n1829), .IN2(n1938), .Q(n280) );
  AND2X1 U3953 ( .IN1(n1842), .IN2(n1865), .Q(n208) );
  AND2X1 U3954 ( .IN1(n1842), .IN2(n1938), .Q(n232) );
  AND2X1 U3957 ( .IN1(n1860), .IN2(n1865), .Q(n64) );
  AND2X1 U3958 ( .IN1(n1860), .IN2(n1938), .Q(n88) );
  AND2X1 U3959 ( .IN1(n1832), .IN2(n1862), .Q(n22) );
  AND2X1 U3960 ( .IN1(n1938), .IN2(n1862), .Q(n40) );
  AND2X1 U3961 ( .IN1(n1915), .IN2(n1865), .Q(n544) );
  AND2X1 U3965 ( .IN1(n1915), .IN2(n1938), .Q(n568) );
  AND2X1 U3966 ( .IN1(n1918), .IN2(n1865), .Q(n496) );
  AND2X1 U3967 ( .IN1(n1918), .IN2(n1938), .Q(n520) );
  AND2X1 U3968 ( .IN1(n1873), .IN2(n1865), .Q(n736) );
  AND2X1 U3971 ( .IN1(n1873), .IN2(n1938), .Q(n760) );
  AND2X1 U3972 ( .IN1(n1898), .IN2(n1865), .Q(n688) );
  AND2X1 U3973 ( .IN1(n1898), .IN2(n1938), .Q(n712) );
  AND2X1 U3974 ( .IN1(n1886), .IN2(n1865), .Q(n640) );
  AND2X1 U3975 ( .IN1(n1886), .IN2(n1938), .Q(n664) );
  AND2X1 U3978 ( .IN1(n1889), .IN2(n1865), .Q(n592) );
  AND2X1 U3979 ( .IN1(n1889), .IN2(n1938), .Q(n616) );
  AND2X1 U3980 ( .IN1(n1905), .IN2(n1865), .Q(n448) );
  AND2X1 U3981 ( .IN1(n1905), .IN2(n1938), .Q(n472) );
  AND2X1 U3982 ( .IN1(n1908), .IN2(n1865), .Q(n400) );
  AND2X1 U3985 ( .IN1(n1908), .IN2(n1938), .Q(n424) );
  AND2X1 U3986 ( .IN1(n1924), .IN2(n1961), .Q(n1936) );
  AND2X1 U3987 ( .IN1(n1924), .IN2(n1962), .Q(n1832) );
  AND2X1 U3988 ( .IN1(n1920), .IN2(n1921), .Q(n1835) );
  AND2X1 U3989 ( .IN1(n1920), .IN2(n1924), .Q(n1841) );
  AND2X1 U3990 ( .IN1(n1920), .IN2(n1925), .Q(n1838) );
  AND2X1 U3994 ( .IN1(n1920), .IN2(n1923), .Q(n1939) );
  AND2X1 U3995 ( .IN1(n1922), .IN2(n1923), .Q(n1836) );
  AND2X1 U3996 ( .IN1(n1923), .IN2(n1962), .Q(n1831) );
  AND2X1 U3997 ( .IN1(n1961), .IN2(n1921), .Q(n1830) );
  AND2X1 U4000 ( .IN1(n1925), .IN2(n1961), .Q(n1833) );
  AND2X1 U4001 ( .IN1(n1922), .IN2(n1921), .Q(n1937) );
  AND2X1 U4002 ( .IN1(n1922), .IN2(n1924), .Q(n1837) );
  AND2X1 U4003 ( .IN1(n1923), .IN2(n1961), .Q(n1866) );
  AND2X1 U4006 ( .IN1(n1925), .IN2(n1962), .Q(n1865) );
  AND2X1 U4007 ( .IN1(n1922), .IN2(n1925), .Q(n1938) );
  AND2X1 U4008 ( .IN1(n1971), .IN2(n1964), .Q(n1840) );
  AND2X1 U4009 ( .IN1(n1988), .IN2(n1951), .Q(n1886) );
  AND2X1 U4010 ( .IN1(n1988), .IN2(n1971), .Q(n1873) );
  AND2X1 U4011 ( .IN1(n1988), .IN2(n1953), .Q(n1898) );
  AND2X1 U4012 ( .IN1(n1988), .IN2(n1943), .Q(n1889) );
  AND2X1 U4015 ( .IN1(n1951), .IN2(n1964), .Q(n1860) );
  AND2X1 U4016 ( .IN1(n1953), .IN2(n1964), .Q(n1861) );
  AND2X1 U4017 ( .IN1(n1942), .IN2(n1951), .Q(n1829) );
  AND2X1 U4018 ( .IN1(n1942), .IN2(n1971), .Q(n1850) );
  AND2X1 U4019 ( .IN1(n1942), .IN2(n1953), .Q(n1853) );
  AND2X1 U4020 ( .IN1(n1942), .IN2(n1943), .Q(n1842) );
  AND2X1 U4024 ( .IN1(n2005), .IN2(n1951), .Q(n1905) );
  AND2X1 U4025 ( .IN1(n2005), .IN2(n1971), .Q(n1915) );
  AND2X1 U4026 ( .IN1(n2005), .IN2(n1953), .Q(n1918) );
  AND2X1 U4027 ( .IN1(n2005), .IN2(n1943), .Q(n1908) );
  NOR2X0 U4030 ( .IN1(n4168), .IN2(n4167), .QN(n1921) );
  NOR2X0 U4031 ( .IN1(n4171), .IN2(n4170), .QN(n1943) );
  NOR2X0 U4032 ( .IN1(n4169), .IN2(n684), .QN(n1962) );
  NOR2X0 U4033 ( .IN1(n4173), .IN2(n4172), .QN(n1964) );
  NOR4X0 U4034 ( .IN1(n813), .IN2(n814), .IN3(n815), .IN4(n816), .QN(n775) );
  NOR4X0 U4035 ( .IN1(n962), .IN2(n963), .IN3(n964), .IN4(n965), .QN(n924) );
  NOR4X0 U4038 ( .IN1(n1111), .IN2(n1112), .IN3(n1113), .IN4(n1114), .QN(n1073) );
  NOR4X0 U4039 ( .IN1(n1260), .IN2(n1261), .IN3(n1262), .IN4(n1263), .QN(n1222) );
  NOR4X0 U4040 ( .IN1(n1409), .IN2(n1410), .IN3(n1411), .IN4(n1412), .QN(n1371) );
  NOR4X0 U4041 ( .IN1(n1558), .IN2(n1559), .IN3(n1560), .IN4(n1561), .QN(n1520) );
  NOR4X0 U4042 ( .IN1(n1707), .IN2(n1708), .IN3(n1709), .IN4(n1710), .QN(n1669) );
  NOR4X0 U4043 ( .IN1(n1877), .IN2(n1878), .IN3(n1879), .IN4(n1880), .QN(n1818) );
  NOR4X0 U4044 ( .IN1(n777), .IN2(n778), .IN3(n779), .IN4(n780), .QN(n776) );
  NOR4X0 U4045 ( .IN1(n926), .IN2(n927), .IN3(n928), .IN4(n929), .QN(n925) );
  NOR4X0 U4046 ( .IN1(n1075), .IN2(n1076), .IN3(n1077), .IN4(n1078), .QN(n1074) );
  NOR4X0 U4047 ( .IN1(n1224), .IN2(n1225), .IN3(n1226), .IN4(n1227), .QN(n1223) );
  NOR4X0 U4048 ( .IN1(n1373), .IN2(n1374), .IN3(n1375), .IN4(n1376), .QN(n1372) );
  NOR4X0 U4049 ( .IN1(n1522), .IN2(n1523), .IN3(n1524), .IN4(n1525), .QN(n1521) );
  NOR4X0 U4052 ( .IN1(n1671), .IN2(n1672), .IN3(n1673), .IN4(n1674), .QN(n1670) );
  NOR4X0 U4053 ( .IN1(n1820), .IN2(n1821), .IN3(n1822), .IN4(n1823), .QN(n1819) );
  INVX0 U4054 ( .IN(n66), .QN(n63) );
  INVX0 U4055 ( .IN(n99), .QN(n96) );
  INVX0 U4056 ( .IN(n132), .QN(n129) );
  INVX0 U4057 ( .IN(n165), .QN(n162) );
  INVX0 U4058 ( .IN(n198), .QN(n195) );
  INVX0 U4059 ( .IN(n231), .QN(n228) );
  INVX0 U4060 ( .IN(n264), .QN(n261) );
  INVX0 U4061 ( .IN(n297), .QN(n294) );
  INVX0 U4062 ( .IN(n66), .QN(n60) );
  INVX0 U4063 ( .IN(n99), .QN(n93) );
  INVX0 U4064 ( .IN(n132), .QN(n126) );
  INVX0 U4065 ( .IN(n165), .QN(n159) );
  INVX0 U4066 ( .IN(n198), .QN(n192) );
  INVX0 U4067 ( .IN(n231), .QN(n225) );
  INVX0 U4068 ( .IN(n264), .QN(n258) );
  INVX0 U4069 ( .IN(n297), .QN(n291) );
  INVX0 U4070 ( .IN(n66), .QN(n57) );
  INVX0 U4071 ( .IN(n99), .QN(n90) );
  INVX0 U4072 ( .IN(n132), .QN(n123) );
  INVX0 U4073 ( .IN(n165), .QN(n156) );
  INVX0 U4074 ( .IN(n198), .QN(n189) );
  INVX0 U4075 ( .IN(n231), .QN(n222) );
  INVX0 U4076 ( .IN(n264), .QN(n255) );
  INVX0 U4077 ( .IN(n297), .QN(n288) );
  INVX0 U4078 ( .IN(n66), .QN(n54) );
  INVX0 U4079 ( .IN(n99), .QN(n87) );
  INVX0 U4080 ( .IN(n132), .QN(n120) );
  INVX0 U4081 ( .IN(n165), .QN(n153) );
  INVX0 U4082 ( .IN(n198), .QN(n186) );
  INVX0 U4083 ( .IN(n231), .QN(n219) );
  INVX0 U4084 ( .IN(n264), .QN(n252) );
  INVX0 U4085 ( .IN(n297), .QN(n285) );
  INVX0 U4086 ( .IN(n66), .QN(n51) );
  INVX0 U4087 ( .IN(n99), .QN(n84) );
  INVX0 U4088 ( .IN(n132), .QN(n117) );
  INVX0 U4089 ( .IN(n165), .QN(n150) );
  INVX0 U4090 ( .IN(n198), .QN(n183) );
  INVX0 U4091 ( .IN(n231), .QN(n216) );
  INVX0 U4092 ( .IN(n264), .QN(n249) );
  INVX0 U4093 ( .IN(n297), .QN(n282) );
  INVX0 U4094 ( .IN(n66), .QN(n48) );
  INVX0 U4095 ( .IN(n99), .QN(n81) );
  INVX0 U4096 ( .IN(n132), .QN(n114) );
  INVX0 U4097 ( .IN(n165), .QN(n147) );
  INVX0 U4098 ( .IN(n198), .QN(n180) );
  INVX0 U4099 ( .IN(n231), .QN(n213) );
  INVX0 U4100 ( .IN(n264), .QN(n246) );
  INVX0 U4101 ( .IN(n297), .QN(n279) );
  INVX0 U4102 ( .IN(n66), .QN(n45) );
  INVX0 U4103 ( .IN(n99), .QN(n78) );
  INVX0 U4104 ( .IN(n132), .QN(n111) );
  INVX0 U4105 ( .IN(n165), .QN(n144) );
  INVX0 U4106 ( .IN(n198), .QN(n177) );
  INVX0 U4107 ( .IN(n231), .QN(n210) );
  INVX0 U4108 ( .IN(n264), .QN(n243) );
  INVX0 U4109 ( .IN(n297), .QN(n276) );
  INVX0 U4110 ( .IN(n66), .QN(n42) );
  INVX0 U4111 ( .IN(n99), .QN(n75) );
  INVX0 U4112 ( .IN(n132), .QN(n108) );
  INVX0 U4113 ( .IN(n165), .QN(n141) );
  INVX0 U4114 ( .IN(n198), .QN(n174) );
  INVX0 U4115 ( .IN(n231), .QN(n207) );
  INVX0 U4116 ( .IN(n264), .QN(n240) );
  INVX0 U4117 ( .IN(n297), .QN(n273) );
  INVX0 U4118 ( .IN(n66), .QN(n39) );
  INVX0 U4119 ( .IN(n99), .QN(n72) );
  INVX0 U4120 ( .IN(n132), .QN(n105) );
  INVX0 U4121 ( .IN(n165), .QN(n138) );
  INVX0 U4122 ( .IN(n198), .QN(n171) );
  INVX0 U4123 ( .IN(n231), .QN(n204) );
  INVX0 U4124 ( .IN(n264), .QN(n237) );
  INVX0 U4125 ( .IN(n297), .QN(n270) );
  INVX0 U4126 ( .IN(n66), .QN(n36) );
  INVX0 U4127 ( .IN(n99), .QN(n69) );
  INVX0 U4128 ( .IN(n132), .QN(n102) );
  INVX0 U4129 ( .IN(n165), .QN(n135) );
  INVX0 U4130 ( .IN(n198), .QN(n168) );
  INVX0 U4131 ( .IN(n231), .QN(n201) );
  INVX0 U4132 ( .IN(n264), .QN(n234) );
  INVX0 U4133 ( .IN(n297), .QN(n267) );
  NOR2X0 U4134 ( .IN1(address[4]), .IN2(address[5]), .QN(n1971) );
  NOR2X0 U4135 ( .IN1(address[1]), .IN2(address[2]), .QN(n1924) );
  NOR2X0 U4136 ( .IN1(address[0]), .IN2(address[3]), .QN(n1920) );
  NOR2X0 U4137 ( .IN1(address[6]), .IN2(address[7]), .QN(n1988) );
  NOR2X0 U4138 ( .IN1(n4170), .IN2(address[5]), .QN(n1953) );
  NOR2X0 U4139 ( .IN1(n4171), .IN2(address[4]), .QN(n1951) );
  NOR2X0 U4140 ( .IN1(n4169), .IN2(address[0]), .QN(n1961) );
  NOR2X0 U4141 ( .IN1(n4167), .IN2(address[2]), .QN(n1925) );
  NOR2X0 U4142 ( .IN1(n4168), .IN2(address[1]), .QN(n1923) );
  NOR2X0 U4143 ( .IN1(n684), .IN2(address[3]), .QN(n1922) );
  NOR2X0 U4144 ( .IN1(n4173), .IN2(address[6]), .QN(n1942) );
  NOR2X0 U4145 ( .IN1(n4172), .IN2(address[7]), .QN(n2005) );
  INVX0 U4146 ( .IN(address[1]), .QN(n4167) );
  INVX0 U4147 ( .IN(address[0]), .QN(n684) );
  INVX0 U4148 ( .IN(address[4]), .QN(n4170) );
  INVX0 U4149 ( .IN(address[6]), .QN(n4172) );
  INVX0 U4150 ( .IN(address[5]), .QN(n4171) );
  INVX0 U4151 ( .IN(address[2]), .QN(n4168) );
  INVX0 U4152 ( .IN(address[3]), .QN(n4169) );
  INVX0 U4153 ( .IN(address[7]), .QN(n4173) );
  NOR4X0 U4154 ( .IN1(n885), .IN2(n886), .IN3(n887), .IN4(n888), .QN(n773) );
  NOR4X0 U4155 ( .IN1(n849), .IN2(n850), .IN3(n851), .IN4(n852), .QN(n774) );
  NOR4X0 U4156 ( .IN1(n1034), .IN2(n1035), .IN3(n1036), .IN4(n1037), .QN(n922)
         );
  NOR4X0 U4157 ( .IN1(n998), .IN2(n999), .IN3(n1000), .IN4(n1001), .QN(n923)
         );
  NOR4X0 U4158 ( .IN1(n1183), .IN2(n1184), .IN3(n1185), .IN4(n1186), .QN(n1071) );
  NOR4X0 U4159 ( .IN1(n1147), .IN2(n1148), .IN3(n1149), .IN4(n1150), .QN(n1072) );
  NOR4X0 U4160 ( .IN1(n1332), .IN2(n1333), .IN3(n1334), .IN4(n1335), .QN(n1220) );
  NOR4X0 U4161 ( .IN1(n1296), .IN2(n1297), .IN3(n1298), .IN4(n1299), .QN(n1221) );
  NOR4X0 U4162 ( .IN1(n1481), .IN2(n1482), .IN3(n1483), .IN4(n1484), .QN(n1369) );
  NOR4X0 U4163 ( .IN1(n1445), .IN2(n1446), .IN3(n1447), .IN4(n1448), .QN(n1370) );
  NOR4X0 U4164 ( .IN1(n1630), .IN2(n1631), .IN3(n1632), .IN4(n1633), .QN(n1518) );
  NOR4X0 U4165 ( .IN1(n1594), .IN2(n1595), .IN3(n1596), .IN4(n1597), .QN(n1519) );
  NOR4X0 U4166 ( .IN1(n1779), .IN2(n1780), .IN3(n1781), .IN4(n1782), .QN(n1667) );
  NOR4X0 U4167 ( .IN1(n1743), .IN2(n1744), .IN3(n1745), .IN4(n1746), .QN(n1668) );
  NOR4X0 U4168 ( .IN1(n1976), .IN2(n1977), .IN3(n1978), .IN4(n1979), .QN(n1816) );
  NOR4X0 U4169 ( .IN1(n1926), .IN2(n1927), .IN3(n1928), .IN4(n1929), .QN(n1817) );
  INVX0 U4170 ( .IN(datain[0]), .QN(n66) );
  INVX0 U4171 ( .IN(datain[1]), .QN(n99) );
  INVX0 U4172 ( .IN(datain[2]), .QN(n132) );
  INVX0 U4173 ( .IN(datain[3]), .QN(n165) );
  INVX0 U4174 ( .IN(datain[4]), .QN(n198) );
  INVX0 U4175 ( .IN(datain[5]), .QN(n231) );
  INVX0 U4176 ( .IN(datain[6]), .QN(n264) );
  INVX0 U4177 ( .IN(datain[7]), .QN(n297) );
endmodule


module memory_access_1 ( mem_in, clk, mem_out, MEM_RD, MEM_data, MEM_acc_mode, 
        stall_Rd, valid, ret_Mem );
  input [31:0] mem_in;
  output [31:0] mem_out;
  output [1:0] MEM_RD;
  output [7:0] MEM_data;
  output [2:0] MEM_acc_mode;
  output [1:0] stall_Rd;
  input clk;
  output valid, ret_Mem;
  wire   \mem_in[23] , \mem_in[22] , \mem_in[21] , \mem_out[19] ,
         \mem_out[18] , \mem_out[17] , \mem_out[16] , N9, N10, n19, n20, n22,
         n23, n24, n25, n26, \sub_72_aco/carry[6] , \sub_72_aco/carry[5] ,
         \sub_72_aco/carry[4] , \sub_72_aco/carry[3] , \sub_72_aco/carry[2] ,
         \sub_72_aco/carry[1] , \sub_72_aco/B[0] , n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n16, n17, n18, \mem_out[20] , n27;
  wire   [7:0] temp_mem_out;
  assign mem_out[24] = 1'b0;
  assign mem_out[25] = 1'b0;
  assign mem_out[26] = 1'b0;
  assign mem_out[27] = 1'b0;
  assign mem_out[28] = 1'b0;
  assign mem_out[29] = 1'b0;
  assign mem_out[30] = 1'b0;
  assign mem_out[31] = 1'b0;
  assign mem_out[23] = \mem_in[23] ;
  assign \mem_in[23]  = mem_in[23];
  assign ret_Mem = \mem_in[22] ;
  assign mem_out[22] = \mem_in[22] ;
  assign \mem_in[22]  = mem_in[22];
  assign mem_out[21] = \mem_in[21] ;
  assign \mem_in[21]  = mem_in[21];
  assign MEM_acc_mode[1] = \mem_out[19] ;
  assign mem_out[19] = \mem_out[19] ;
  assign MEM_acc_mode[0] = \mem_out[18] ;
  assign mem_out[18] = \mem_out[18] ;
  assign stall_Rd[1] = \mem_out[17] ;
  assign mem_out[17] = \mem_out[17] ;
  assign stall_Rd[0] = \mem_out[16] ;
  assign mem_out[16] = \mem_out[16] ;
  assign MEM_acc_mode[2] = \mem_out[20] ;
  assign mem_out[20] = \mem_out[20] ;

  AND2X1 U42 ( .IN1(temp_mem_out[1]), .IN2(N9), .Q(mem_out[9]) );
  AND2X1 U43 ( .IN1(temp_mem_out[0]), .IN2(N9), .Q(mem_out[8]) );
  AND2X1 U46 ( .IN1(temp_mem_out[7]), .IN2(N9), .Q(mem_out[15]) );
  AND2X1 U47 ( .IN1(temp_mem_out[6]), .IN2(N9), .Q(mem_out[14]) );
  AND2X1 U48 ( .IN1(temp_mem_out[5]), .IN2(N9), .Q(mem_out[13]) );
  AND2X1 U49 ( .IN1(temp_mem_out[4]), .IN2(N9), .Q(mem_out[12]) );
  AND2X1 U50 ( .IN1(temp_mem_out[3]), .IN2(N9), .Q(mem_out[11]) );
  AND2X1 U51 ( .IN1(temp_mem_out[2]), .IN2(N9), .Q(mem_out[10]) );
  AO21X1 U54 ( .IN1(n23), .IN2(mem_in[17]), .IN3(n22), .Q(MEM_RD[1]) );
  AO21X1 U55 ( .IN1(n23), .IN2(mem_in[16]), .IN3(n22), .Q(MEM_RD[0]) );
  AOI21X1 U58 ( .IN1(n24), .IN2(n26), .IN3(mem_in[18]), .QN(n23) );
  data_ram_1 mem_acc ( .clk(clk), .R(N9), .W(N10), .address(mem_in[7:0]), 
        .datain(mem_in[15:8]), .dataout(temp_mem_out) );
  INVX0 U2 ( .IN(mem_in[6]), .QN(n12) );
  INVX0 U3 ( .IN(\mem_in[21] ), .QN(n27) );
  AND2X1 U4 ( .IN1(\mem_out[18] ), .IN2(n18), .Q(N9) );
  AND2X1 U5 ( .IN1(mem_in[16]), .IN2(\mem_in[21] ), .Q(\mem_out[16] ) );
  AND2X1 U6 ( .IN1(mem_in[17]), .IN2(\mem_in[21] ), .Q(\mem_out[17] ) );
  INVX0 U7 ( .IN(n24), .QN(\mem_out[20] ) );
  XOR2X1 U8 ( .IN1(mem_in[7]), .IN2(n9), .Q(n1) );
  XOR2X1 U9 ( .IN1(\sub_72_aco/carry[6] ), .IN2(mem_in[6]), .Q(n2) );
  XOR2X1 U10 ( .IN1(\sub_72_aco/carry[1] ), .IN2(mem_in[1]), .Q(n3) );
  XOR2X1 U11 ( .IN1(\sub_72_aco/carry[5] ), .IN2(mem_in[5]), .Q(n4) );
  XOR2X1 U12 ( .IN1(\sub_72_aco/carry[4] ), .IN2(mem_in[4]), .Q(n5) );
  XOR2X1 U13 ( .IN1(\sub_72_aco/carry[3] ), .IN2(mem_in[3]), .Q(n6) );
  XOR2X1 U14 ( .IN1(\sub_72_aco/carry[2] ), .IN2(mem_in[2]), .Q(n7) );
  XOR2X1 U15 ( .IN1(n20), .IN2(mem_in[0]), .Q(n8) );
  NAND4X0 U16 ( .IN1(mem_in[20]), .IN2(\mem_in[21] ), .IN3(n16), .IN4(n17), 
        .QN(n20) );
  NOR2X0 U17 ( .IN1(n22), .IN2(n23), .QN(n19) );
  NAND2X0 U18 ( .IN1(n11), .IN2(n12), .QN(n9) );
  OR2X1 U19 ( .IN1(\sub_72_aco/B[0] ), .IN2(n10), .Q(N10) );
  AND3X1 U20 ( .IN1(n16), .IN2(n18), .IN3(\mem_out[19] ), .Q(n10) );
  INVX0 U21 ( .IN(n13), .QN(\sub_72_aco/B[0] ) );
  INVX0 U22 ( .IN(\sub_72_aco/carry[6] ), .QN(n11) );
  NAND4X0 U23 ( .IN1(mem_in[19]), .IN2(mem_in[18]), .IN3(\mem_in[21] ), .IN4(
        n18), .QN(n25) );
  INVX0 U24 ( .IN(mem_in[20]), .QN(n18) );
  OR2X1 U25 ( .IN1(\sub_72_aco/carry[2] ), .IN2(mem_in[2]), .Q(
        \sub_72_aco/carry[3] ) );
  OR2X1 U26 ( .IN1(\sub_72_aco/carry[3] ), .IN2(mem_in[3]), .Q(
        \sub_72_aco/carry[4] ) );
  OR2X1 U27 ( .IN1(\sub_72_aco/carry[5] ), .IN2(mem_in[5]), .Q(
        \sub_72_aco/carry[6] ) );
  OR2X1 U28 ( .IN1(n20), .IN2(mem_in[0]), .Q(\sub_72_aco/carry[1] ) );
  OR2X1 U29 ( .IN1(\sub_72_aco/carry[1] ), .IN2(mem_in[1]), .Q(
        \sub_72_aco/carry[2] ) );
  OR2X1 U30 ( .IN1(\sub_72_aco/carry[4] ), .IN2(mem_in[4]), .Q(
        \sub_72_aco/carry[5] ) );
  NAND4X0 U31 ( .IN1(mem_in[20]), .IN2(\mem_in[21] ), .IN3(n16), .IN4(n17), 
        .QN(n13) );
  NOR2X0 U32 ( .IN1(n27), .IN2(n6), .QN(mem_out[3]) );
  NOR2X0 U33 ( .IN1(n27), .IN2(n5), .QN(mem_out[4]) );
  NOR2X0 U34 ( .IN1(n27), .IN2(n4), .QN(mem_out[5]) );
  NOR2X0 U35 ( .IN1(n27), .IN2(n7), .QN(mem_out[2]) );
  NOR2X0 U36 ( .IN1(n27), .IN2(n3), .QN(mem_out[1]) );
  NOR2X0 U37 ( .IN1(n27), .IN2(n2), .QN(mem_out[6]) );
  NOR2X0 U38 ( .IN1(n27), .IN2(n8), .QN(mem_out[0]) );
  NAND2X0 U39 ( .IN1(n25), .IN2(n13), .QN(n22) );
  NOR2X0 U40 ( .IN1(n19), .IN2(n2), .QN(MEM_data[6]) );
  NOR2X0 U41 ( .IN1(n19), .IN2(n4), .QN(MEM_data[5]) );
  NOR2X0 U44 ( .IN1(n19), .IN2(n5), .QN(MEM_data[4]) );
  NOR2X0 U45 ( .IN1(n19), .IN2(n6), .QN(MEM_data[3]) );
  NOR2X0 U52 ( .IN1(n19), .IN2(n7), .QN(MEM_data[2]) );
  NOR2X0 U53 ( .IN1(n19), .IN2(n3), .QN(MEM_data[1]) );
  NOR2X0 U56 ( .IN1(n19), .IN2(n8), .QN(MEM_data[0]) );
  INVX0 U57 ( .IN(n19), .QN(valid) );
  NAND2X0 U59 ( .IN1(mem_in[20]), .IN2(\mem_in[21] ), .QN(n24) );
  NOR2X0 U60 ( .IN1(n27), .IN2(n1), .QN(mem_out[7]) );
  INVX0 U61 ( .IN(mem_in[19]), .QN(n14) );
  NOR2X0 U62 ( .IN1(n17), .IN2(n27), .QN(\mem_out[19] ) );
  INVX0 U63 ( .IN(mem_in[19]), .QN(n17) );
  NAND2X0 U64 ( .IN1(\mem_in[21] ), .IN2(n14), .QN(n26) );
  NOR2X0 U65 ( .IN1(n16), .IN2(n27), .QN(\mem_out[18] ) );
  INVX0 U66 ( .IN(mem_in[18]), .QN(n16) );
  NOR2X0 U67 ( .IN1(n19), .IN2(n1), .QN(MEM_data[7]) );
endmodule


module my_DFF_1_64 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_63 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_62 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_61 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_60 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_59 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_58 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_57 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_56 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_55 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_54 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_53 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_52 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_51 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_50 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_49 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_48 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_47 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_46 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_45 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_44 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_43 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U2 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U3 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_42 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_41 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_40 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_39 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_38 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_37 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_36 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_35 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_34 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_DFF_1_33 ( d, clk, rst, e, q );
  input d, clk, rst, e;
  output q;
  wire   n1, n2, n4;

  DFFARX1 q_reg ( .D(n4), .CLK(clk), .RSTB(n1), .Q(q) );
  AO22X1 U3 ( .IN1(q), .IN2(n2), .IN3(e), .IN4(d), .Q(n4) );
  INVX0 U2 ( .IN(rst), .QN(n1) );
  INVX0 U4 ( .IN(e), .QN(n2) );
endmodule


module my_nDFF_n32_1 ( clk, rst, e, d, q );
  input [31:0] d;
  output [31:0] q;
  input clk, rst, e;
  wire   n1, n2, n3;

  my_DFF_1_64 fx_0 ( .d(d[0]), .clk(clk), .rst(n3), .e(e), .q(q[0]) );
  my_DFF_1_63 fx_1 ( .d(d[1]), .clk(clk), .rst(n3), .e(e), .q(q[1]) );
  my_DFF_1_62 fx_2 ( .d(d[2]), .clk(clk), .rst(n3), .e(e), .q(q[2]) );
  my_DFF_1_61 fx_3 ( .d(d[3]), .clk(clk), .rst(n3), .e(e), .q(q[3]) );
  my_DFF_1_60 fx_4 ( .d(d[4]), .clk(clk), .rst(n3), .e(e), .q(q[4]) );
  my_DFF_1_59 fx_5 ( .d(d[5]), .clk(clk), .rst(n3), .e(e), .q(q[5]) );
  my_DFF_1_58 fx_6 ( .d(d[6]), .clk(clk), .rst(n3), .e(e), .q(q[6]) );
  my_DFF_1_57 fx_7 ( .d(d[7]), .clk(clk), .rst(n3), .e(e), .q(q[7]) );
  my_DFF_1_56 fx_8 ( .d(d[8]), .clk(clk), .rst(n2), .e(e), .q(q[8]) );
  my_DFF_1_55 fx_9 ( .d(d[9]), .clk(clk), .rst(n2), .e(e), .q(q[9]) );
  my_DFF_1_54 fx_10 ( .d(d[10]), .clk(clk), .rst(n2), .e(e), .q(q[10]) );
  my_DFF_1_53 fx_11 ( .d(d[11]), .clk(clk), .rst(n2), .e(e), .q(q[11]) );
  my_DFF_1_52 fx_12 ( .d(d[12]), .clk(clk), .rst(n2), .e(e), .q(q[12]) );
  my_DFF_1_51 fx_13 ( .d(d[13]), .clk(clk), .rst(n2), .e(e), .q(q[13]) );
  my_DFF_1_50 fx_14 ( .d(d[14]), .clk(clk), .rst(n2), .e(e), .q(q[14]) );
  my_DFF_1_49 fx_15 ( .d(d[15]), .clk(clk), .rst(n2), .e(e), .q(q[15]) );
  my_DFF_1_48 fx_16 ( .d(d[16]), .clk(clk), .rst(n2), .e(e), .q(q[16]) );
  my_DFF_1_47 fx_17 ( .d(d[17]), .clk(clk), .rst(n2), .e(e), .q(q[17]) );
  my_DFF_1_46 fx_18 ( .d(d[18]), .clk(clk), .rst(n2), .e(e), .q(q[18]) );
  my_DFF_1_45 fx_19 ( .d(d[19]), .clk(clk), .rst(n2), .e(e), .q(q[19]) );
  my_DFF_1_44 fx_20 ( .d(d[20]), .clk(clk), .rst(n1), .e(e), .q(q[20]) );
  my_DFF_1_43 fx_21 ( .d(d[21]), .clk(clk), .rst(n1), .e(e), .q(q[21]) );
  my_DFF_1_42 fx_22 ( .d(d[22]), .clk(clk), .rst(n1), .e(e), .q(q[22]) );
  my_DFF_1_41 fx_23 ( .d(d[23]), .clk(clk), .rst(n1), .e(e), .q(q[23]) );
  my_DFF_1_40 fx_24 ( .d(d[24]), .clk(clk), .rst(n1), .e(e), .q(q[24]) );
  my_DFF_1_39 fx_25 ( .d(d[25]), .clk(clk), .rst(n1), .e(e), .q(q[25]) );
  my_DFF_1_38 fx_26 ( .d(d[26]), .clk(clk), .rst(n1), .e(e), .q(q[26]) );
  my_DFF_1_37 fx_27 ( .d(d[27]), .clk(clk), .rst(n1), .e(e), .q(q[27]) );
  my_DFF_1_36 fx_28 ( .d(d[28]), .clk(clk), .rst(n1), .e(e), .q(q[28]) );
  my_DFF_1_35 fx_29 ( .d(d[29]), .clk(clk), .rst(n1), .e(e), .q(q[29]) );
  my_DFF_1_34 fx_30 ( .d(d[30]), .clk(clk), .rst(n1), .e(e), .q(q[30]) );
  my_DFF_1_33 fx_31 ( .d(d[31]), .clk(clk), .rst(n1), .e(e), .q(q[31]) );
  NBUFFX2 U1 ( .IN(rst), .Q(n2) );
  NBUFFX2 U2 ( .IN(rst), .Q(n1) );
  NBUFFX2 U3 ( .IN(rst), .Q(n3) );
endmodule


module write_back_1 ( write_in, clk, W, SP_EN, Rd, data, SP_in, port_out, 
        valid, ret_WB, pop_flags );
  input [31:0] write_in;
  output [1:0] Rd;
  output [7:0] data;
  output [7:0] SP_in;
  output [7:0] port_out;
  input clk;
  output W, SP_EN, valid, ret_WB, pop_flags;
  wire   write_in_23, write_in_22, write_in_21, write_in_20, write_in_19,
         write_in_18, \write_in[17] , \write_in[16] , N4, N18, N19, n6, n7, n8,
         n9, n10, n11, n12, n13, n1, n2, n3, n4, n5;
  assign pop_flags = write_in_23;
  assign write_in_23 = write_in[23];
  assign ret_WB = write_in_22;
  assign write_in_22 = write_in[22];
  assign write_in_21 = write_in[21];
  assign write_in_20 = write_in[20];
  assign write_in_19 = write_in[19];
  assign write_in_18 = write_in[18];
  assign Rd[1] = \write_in[17] ;
  assign \write_in[17]  = write_in[17];
  assign Rd[0] = \write_in[16] ;
  assign \write_in[16]  = write_in[16];
  assign SP_EN = N4;
  assign W = N19;

  LATCHX1 \temp_port_reg[7]  ( .CLK(N18), .D(write_in[7]), .Q(port_out[7]) );
  LATCHX1 \temp_port_reg[6]  ( .CLK(N18), .D(write_in[6]), .Q(port_out[6]) );
  LATCHX1 \temp_port_reg[5]  ( .CLK(N18), .D(write_in[5]), .Q(port_out[5]) );
  LATCHX1 \temp_port_reg[4]  ( .CLK(N18), .D(write_in[4]), .Q(port_out[4]) );
  LATCHX1 \temp_port_reg[3]  ( .CLK(N18), .D(write_in[3]), .Q(port_out[3]) );
  LATCHX1 \temp_port_reg[2]  ( .CLK(N18), .D(write_in[2]), .Q(port_out[2]) );
  LATCHX1 \temp_port_reg[1]  ( .CLK(N18), .D(write_in[1]), .Q(port_out[1]) );
  LATCHX1 \temp_port_reg[0]  ( .CLK(N18), .D(write_in[0]), .Q(port_out[0]) );
  AND3X1 U9 ( .IN1(n6), .IN2(n7), .IN3(write_in_21), .Q(valid) );
  NAND3X0 U10 ( .IN1(n1), .IN2(n4), .IN3(write_in_19), .QN(n6) );
  AO22X1 U11 ( .IN1(write_in[7]), .IN2(n8), .IN3(write_in[15]), .IN4(n2), .Q(
        data[7]) );
  AO22X1 U12 ( .IN1(write_in[6]), .IN2(n8), .IN3(write_in[14]), .IN4(n2), .Q(
        data[6]) );
  AO22X1 U13 ( .IN1(write_in[5]), .IN2(n8), .IN3(write_in[13]), .IN4(n2), .Q(
        data[5]) );
  AO22X1 U14 ( .IN1(write_in[4]), .IN2(n8), .IN3(write_in[12]), .IN4(n2), .Q(
        data[4]) );
  AO22X1 U15 ( .IN1(write_in[3]), .IN2(n8), .IN3(write_in[11]), .IN4(n2), .Q(
        data[3]) );
  AO22X1 U16 ( .IN1(write_in[2]), .IN2(n8), .IN3(write_in[10]), .IN4(n2), .Q(
        data[2]) );
  AO22X1 U17 ( .IN1(write_in[1]), .IN2(n8), .IN3(write_in[9]), .IN4(n2), .Q(
        data[1]) );
  AO22X1 U18 ( .IN1(write_in[0]), .IN2(n8), .IN3(write_in[8]), .IN4(n2), .Q(
        data[0]) );
  AND3X1 U19 ( .IN1(write_in_21), .IN2(n1), .IN3(n10), .Q(n8) );
  XOR2X1 U20 ( .IN1(n3), .IN2(write_in_20), .Q(n10) );
  AND2X1 U21 ( .IN1(N4), .IN2(write_in[7]), .Q(SP_in[7]) );
  AND2X1 U22 ( .IN1(N4), .IN2(write_in[6]), .Q(SP_in[6]) );
  AND2X1 U23 ( .IN1(N4), .IN2(write_in[5]), .Q(SP_in[5]) );
  AND2X1 U24 ( .IN1(N4), .IN2(write_in[4]), .Q(SP_in[4]) );
  AND2X1 U25 ( .IN1(N4), .IN2(write_in[3]), .Q(SP_in[3]) );
  AND2X1 U26 ( .IN1(N4), .IN2(write_in[2]), .Q(SP_in[2]) );
  AND2X1 U27 ( .IN1(N4), .IN2(write_in[1]), .Q(SP_in[1]) );
  AND2X1 U28 ( .IN1(N4), .IN2(write_in[0]), .Q(SP_in[0]) );
  NOR3X0 U30 ( .IN1(n12), .IN2(write_in_23), .IN3(write_in_22), .QN(N19) );
  OA221X1 U31 ( .IN1(n3), .IN2(n11), .IN3(n5), .IN4(n13), .IN5(n9), .Q(n12) );
  NAND3X0 U32 ( .IN1(write_in_18), .IN2(n4), .IN3(write_in_21), .QN(n9) );
  NAND3X0 U33 ( .IN1(write_in_20), .IN2(n1), .IN3(write_in_21), .QN(n11) );
  NOR3X0 U34 ( .IN1(n7), .IN2(write_in_19), .IN3(n5), .QN(N18) );
  INVX0 U2 ( .IN(n9), .QN(n2) );
  INVX0 U3 ( .IN(write_in_19), .QN(n3) );
  INVX0 U4 ( .IN(write_in_20), .QN(n4) );
  INVX0 U5 ( .IN(write_in_18), .QN(n1) );
  NAND2X0 U6 ( .IN1(write_in_20), .IN2(write_in_18), .QN(n7) );
  NAND2X0 U7 ( .IN1(n3), .IN2(n4), .QN(n13) );
  INVX0 U8 ( .IN(write_in_21), .QN(n5) );
  OAI22X2 U29 ( .IN1(n9), .IN2(n3), .IN3(n11), .IN4(write_in_19), .QN(N4) );
endmodule


module CPU ( clk, rst, INT_IN, IN_PORT, OUT_PORT );
  input [7:0] IN_PORT;
  output [7:0] OUT_PORT;
  input clk, rst, INT_IN;
  wire   inst_R, stall_en, stall, ret_Ex, ret_Mem, ret_WB, branch, EX_RTI,
         imm_en, PC_src, return_address_src, flags_src, reg_W, SP_EN,
         ID_EXin_57, ID_EXin_56, ID_EXin_42, ID_EXin_41, ID_EXin_40,
         ID_EXin_39, ID_EXin_38, ID_EXin_34, MEM_valid, WB_valid, pop_flags,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n47, n48, n49, n50;
  wire   [7:0] PCin;
  wire   [25:0] IF_IDin;
  wire   [31:0] IF_ID;
  wire   [7:0] WB_data;
  wire   [7:0] target_address;
  wire   [1:0] Rs1;
  wire   [1:0] Rs2;
  wire   [1:0] Rd;
  wire   [2:0] acc_mode;
  wire   [7:0] offset;
  wire   [3:0] alu_op;
  wire   [2:0] branch_mode;
  wire   [1:0] WB_Rd;
  wire   [7:0] SP_IN;
  wire   [7:0] S1;
  wire   [7:0] S2;
  wire   [17:10] ID_EXin;
  wire   [3:0] flags_input;
  wire   [63:0] ID_EX;
  wire   [3:0] flags;
  wire   [7:0] MEM_data;
  wire   [1:0] MEM_Rd;
  wire   [2:0] MEM_acc_mode;
  wire   [1:0] stall_Rd;
  wire   [31:0] EX_MEMin;
  wire   [3:0] flags_in;
  wire   [31:0] EX_MEM;
  wire   [31:0] MEM_WBin;
  wire   [31:0] MEM_WB;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22;

  AO222X1 U45 ( .IN1(n17), .IN2(PCin[7]), .IN3(S2[7]), .IN4(n18), .IN5(
        return_address_src), .IN6(IF_IDin[25]), .Q(ID_EXin[17]) );
  AO222X1 U46 ( .IN1(n17), .IN2(PCin[6]), .IN3(S2[6]), .IN4(n18), .IN5(
        IF_IDin[24]), .IN6(return_address_src), .Q(ID_EXin[16]) );
  AO222X1 U47 ( .IN1(n17), .IN2(PCin[5]), .IN3(S2[5]), .IN4(n18), .IN5(
        IF_IDin[23]), .IN6(return_address_src), .Q(ID_EXin[15]) );
  AO222X1 U48 ( .IN1(n17), .IN2(PCin[4]), .IN3(S2[4]), .IN4(n18), .IN5(
        IF_IDin[22]), .IN6(return_address_src), .Q(ID_EXin[14]) );
  AO221X1 U49 ( .IN1(n19), .IN2(flags_input[3]), .IN3(S2[3]), .IN4(n18), .IN5(
        n20), .Q(ID_EXin[13]) );
  AO22X1 U50 ( .IN1(IF_IDin[21]), .IN2(return_address_src), .IN3(PCin[3]), 
        .IN4(n17), .Q(n20) );
  AO22X1 U51 ( .IN1(flags_in[3]), .IN2(n50), .IN3(pop_flags), .IN4(WB_data[3]), 
        .Q(flags_input[3]) );
  AO22X1 U54 ( .IN1(flags_in[2]), .IN2(n50), .IN3(WB_data[2]), .IN4(pop_flags), 
        .Q(flags_input[2]) );
  AO221X1 U55 ( .IN1(n19), .IN2(flags_input[1]), .IN3(S2[1]), .IN4(n18), .IN5(
        n22), .Q(ID_EXin[11]) );
  AO22X1 U56 ( .IN1(IF_IDin[19]), .IN2(return_address_src), .IN3(PCin[1]), 
        .IN4(n17), .Q(n22) );
  AO22X1 U57 ( .IN1(flags_in[1]), .IN2(n50), .IN3(WB_data[1]), .IN4(pop_flags), 
        .Q(flags_input[1]) );
  AO221X1 U58 ( .IN1(n19), .IN2(flags_input[0]), .IN3(S2[0]), .IN4(n18), .IN5(
        n23), .Q(ID_EXin[10]) );
  AO22X1 U59 ( .IN1(IF_IDin[18]), .IN2(return_address_src), .IN3(n17), .IN4(
        PCin[0]), .Q(n23) );
  AND2X1 U60 ( .IN1(PC_src), .IN2(n24), .Q(n17) );
  AO22X1 U61 ( .IN1(flags_in[0]), .IN2(n50), .IN3(WB_data[0]), .IN4(pop_flags), 
        .Q(flags_input[0]) );
  my_nDFF_n8_0 PC_reg ( .clk(clk), .rst(rst), .e(1'b1), .d(PCin) );
  inst_ram_1 inst_mem ( .clk(clk), .R(inst_R), .address(PCin) );
  my_nDFF_n32_0 IF_ID_reg ( .clk(clk), .rst(1'b0), .e(stall_en), .d({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, IF_IDin[25:8], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .q(IF_ID) );
  CU CU_comp ( .clk(clk), .rst(rst), .INT_IN(INT_IN), .stall(stall), .ret_Ex(
        ret_Ex), .ret_Mem(ret_Mem), .ret_WB(ret_WB), .branch(branch), .EX_RTI(
        EX_RTI), .ret_PC(WB_data), .target_address(target_address), .IF_ID(
        IF_ID), .inst_R(inst_R), .stall_en(stall_en), .f1_en(ID_EXin_40), 
        .f2_en(ID_EXin_41), .imm_en(imm_en), .Rs1(Rs1), .Rs2(Rs2), .Rd(Rd), 
        .acc_mode(acc_mode), .NOP(ID_EXin_38), .offset_en(ID_EXin_34), 
        .offset({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, offset[0]}), .alu_op(alu_op), .change_flags(
        ID_EXin_39), .branch_mode(branch_mode), .ret(ID_EXin_42), .PC_src(
        PC_src), .push_PC(IF_IDin[17]), .push_flags(IF_IDin[16]), 
        .return_address(IF_IDin[25:18]), .return_address_src(
        return_address_src), .flags_src(flags_src), .pre_RTI(ID_EXin_56), 
        .pre_pop_flags(ID_EXin_57), .PCin(PCin) );
  reg_file_1 Registers_file ( .clk(clk), .rst(rst), .R(1'b1), .W(reg_W), 
        .SP_EN(SP_EN), .Rs1(Rs1), .Rs2(Rs2), .Rd(WB_Rd), .data_sp(SP_IN), 
        .data(WB_data), .S1(S1), .S2(S2) );
  my_nDFF_n64 ID_EX_reg ( .clk(clk), .rst(rst), .e(stall_en), .d({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, ID_EXin_57, ID_EXin_56, S2, Rs2, branch_mode, 
        ID_EXin_42, ID_EXin_41, ID_EXin_40, ID_EXin_39, ID_EXin_38, acc_mode, 
        ID_EXin_34, Rd, alu_op, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        offset[0], Rs2, ID_EXin, Rs1, n32, n31, n30, n29, n28, n27, n26, n25}), 
        .q(ID_EX) );
  execute_1 Eexecute_unit ( .ID_EX(ID_EX), .flags_in(flags), .mem_data(
        MEM_data), .mem_rd(MEM_Rd), .mem_acc_mode(MEM_acc_mode), .stall_Rd(
        stall_Rd), .mem_valid(MEM_valid), .wb_data(WB_data), .wb_rd(WB_Rd), 
        .wb_valid(WB_valid), .sp_data(SP_IN), .sp_en(SP_EN), .IN_PORT(IN_PORT), 
        .EX_MEM({SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, EX_MEMin[23:0]}), 
        .flags_out(flags_in), .stall(stall), .ret_ex(ret_Ex), .branch(branch), 
        .target_addr(target_address), .rti(EX_RTI) );
  my_nDFF_n4 flags_reg ( .clk(clk), .rst(rst), .e(1'b1), .d(flags_input), .q(
        flags) );
  my_nDFF_n32_2 EX_MEM_reg ( .clk(clk), .rst(rst), .e(1'b1), .d({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, EX_MEMin[23:0]}), .q(EX_MEM) );
  memory_access_1 memory_access_unit ( .mem_in(EX_MEM), .clk(clk), .mem_out({
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, MEM_WBin[23:0]}), 
        .MEM_RD(MEM_Rd), .MEM_data(MEM_data), .MEM_acc_mode(MEM_acc_mode), 
        .stall_Rd(stall_Rd), .valid(MEM_valid), .ret_Mem(ret_Mem) );
  my_nDFF_n32_1 MEM_WB_reg ( .clk(clk), .rst(rst), .e(1'b1), .d({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, MEM_WBin[23:0]}), .q(MEM_WB) );
  write_back_1 write_back_unit ( .write_in(MEM_WB), .clk(clk), .W(reg_W), 
        .SP_EN(SP_EN), .Rd(WB_Rd), .data(WB_data), .SP_in(SP_IN), .port_out(
        OUT_PORT), .valid(WB_valid), .ret_WB(ret_WB), .pop_flags(pop_flags) );
  AND2X1 U62 ( .IN1(S1[0]), .IN2(n47), .Q(n25) );
  AND2X1 U63 ( .IN1(S1[1]), .IN2(n47), .Q(n26) );
  AND2X1 U64 ( .IN1(S1[2]), .IN2(n47), .Q(n27) );
  AND2X1 U65 ( .IN1(S1[3]), .IN2(n47), .Q(n28) );
  AND2X1 U66 ( .IN1(S1[4]), .IN2(n47), .Q(n29) );
  AND2X1 U67 ( .IN1(S1[5]), .IN2(n47), .Q(n30) );
  AND2X1 U68 ( .IN1(S1[6]), .IN2(n47), .Q(n31) );
  AND2X1 U69 ( .IN1(S1[7]), .IN2(n47), .Q(n32) );
  AND2X1 U70 ( .IN1(n19), .IN2(flags_input[2]), .Q(n33) );
  AND2X1 U71 ( .IN1(S2[2]), .IN2(n18), .Q(n34) );
  OR3X1 U72 ( .IN1(n33), .IN2(n34), .IN3(n21), .Q(ID_EXin[12]) );
  INVX0 U73 ( .IN(imm_en), .QN(n47) );
  NOR2X0 U74 ( .IN1(n49), .IN2(PC_src), .QN(n18) );
  INVX0 U75 ( .IN(n24), .QN(n49) );
  NAND2X0 U76 ( .IN1(IF_IDin[20]), .IN2(return_address_src), .QN(n35) );
  NAND2X0 U77 ( .IN1(n37), .IN2(n44), .QN(IF_IDin[9]) );
  NAND2X0 U78 ( .IN1(n37), .IN2(n42), .QN(IF_IDin[11]) );
  INVX0 U79 ( .IN(PCin[3]), .QN(n42) );
  NAND2X0 U80 ( .IN1(n37), .IN2(n43), .QN(IF_IDin[10]) );
  INVX0 U81 ( .IN(PCin[2]), .QN(n43) );
  NAND2X0 U82 ( .IN1(n37), .IN2(n45), .QN(IF_IDin[8]) );
  INVX0 U83 ( .IN(PCin[0]), .QN(n45) );
  NAND2X0 U84 ( .IN1(n37), .IN2(n41), .QN(IF_IDin[12]) );
  INVX0 U85 ( .IN(PCin[4]), .QN(n41) );
  NAND2X0 U86 ( .IN1(n37), .IN2(n40), .QN(IF_IDin[13]) );
  INVX0 U87 ( .IN(PCin[5]), .QN(n40) );
  NAND2X0 U88 ( .IN1(n37), .IN2(n39), .QN(IF_IDin[14]) );
  INVX0 U89 ( .IN(PCin[6]), .QN(n39) );
  NAND2X0 U90 ( .IN1(n37), .IN2(n38), .QN(IF_IDin[15]) );
  INVX0 U91 ( .IN(PCin[7]), .QN(n38) );
  NOR2X0 U92 ( .IN1(n48), .IN2(return_address_src), .QN(n19) );
  INVX0 U93 ( .IN(flags_src), .QN(n48) );
  NOR2X0 U94 ( .IN1(flags_src), .IN2(return_address_src), .QN(n24) );
  INVX0 U95 ( .IN(pop_flags), .QN(n50) );
  INVX0 U96 ( .IN(rst), .QN(n37) );
  NAND2X0 U97 ( .IN1(PCin[2]), .IN2(n17), .QN(n36) );
  NAND2X0 U98 ( .IN1(n35), .IN2(n36), .QN(n21) );
  INVX0 U99 ( .IN(PCin[1]), .QN(n44) );
endmodule

